/afs/ece.cmu.edu/project/km_group/.vol9/asap7/fpga_demos/simple_fpga/mux_BB.lef