module Alu(
  input         clock,
  input         reset,
  input  [15:0] io_i0,
  input  [15:0] io_i1,
  input  [31:0] io_ib32,
  input  [7:0]  io_ctrl,
  output [15:0] io_q,
  output [31:0] io_ob32,
  input  [31:0] io_config,
  input         io_gndOuts,
  input         io_clkEnb
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  _i0FF_T = ~io_clkEnb; // @[CLBlut4N10Alu.scala 97:44]
  reg [15:0] i0FF; // @[Reg.scala 28:20]
  reg [15:0] i1FF; // @[Reg.scala 28:20]
  reg [31:0] ib32FF; // @[Reg.scala 28:20]
  wire [15:0] in0 = io_config[0] ? io_i0 : i0FF; // @[CLBlut4N10Alu.scala 101:16]
  wire [15:0] in1 = io_config[1] ? io_i1 : i1FF; // @[CLBlut4N10Alu.scala 102:16]
  wire [31:0] ib32 = io_config[2] ? io_ib32 : ib32FF; // @[CLBlut4N10Alu.scala 103:17]
  wire [15:0] _acc_T_1 = in0 + in1; // @[CLBlut4N10Alu.scala 105:17]
  wire [31:0] _GEN_4 = {{16'd0}, _acc_T_1}; // @[CLBlut4N10Alu.scala 105:23]
  wire [31:0] acc = _GEN_4 + ib32; // @[CLBlut4N10Alu.scala 105:23]
  wire  _accFF_T_4 = io_ctrl[1] & _i0FF_T; // @[CLBlut4N10Alu.scala 107:68]
  reg [31:0] accFF; // @[Reg.scala 28:20]
  wire [31:0] _out_T_1 = io_config[3] ? accFF : acc; // @[CLBlut4N10Alu.scala 110:16]
  wire  _out_T_2 = ~io_gndOuts; // @[CLBlut4N10Alu.scala 110:45]
  wire [31:0] _GEN_5 = {{31'd0}, _out_T_2}; // @[CLBlut4N10Alu.scala 110:43]
  wire [31:0] out = _out_T_1 & _GEN_5; // @[CLBlut4N10Alu.scala 110:43]
  assign io_q = io_ctrl[1] ? out[31:16] : out[15:0]; // @[CLBlut4N10Alu.scala 112:14]
  assign io_ob32 = _out_T_1 & _GEN_5; // @[CLBlut4N10Alu.scala 110:43]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      i0FF <= 16'h0; // @[Reg.scala 28:20]
    end else if (_i0FF_T) begin // @[Reg.scala 29:18]
      i0FF <= io_i0; // @[Reg.scala 29:22]
    end
    if (reset) begin // @[Reg.scala 28:20]
      i1FF <= 16'h0; // @[Reg.scala 28:20]
    end else if (_i0FF_T) begin // @[Reg.scala 29:18]
      i1FF <= io_i1; // @[Reg.scala 29:22]
    end
    if (reset) begin // @[Reg.scala 28:20]
      ib32FF <= 32'h0; // @[Reg.scala 28:20]
    end else if (_i0FF_T) begin // @[Reg.scala 29:18]
      ib32FF <= io_ib32; // @[Reg.scala 29:22]
    end
    if (reset) begin // @[Reg.scala 28:20]
      accFF <= 32'h0; // @[Reg.scala 28:20]
    end else if (_accFF_T_4) begin // @[Reg.scala 29:18]
      if (io_ctrl[0]) begin // @[CLBlut4N10Alu.scala 107:28]
        accFF <= 32'h0;
      end else begin
        accFF <= acc;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i0FF = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  i1FF = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  ib32FF = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  accFF = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Ble4(
  input         clock,
  input         reset,
  input  [19:0] io_config,
  input         io_in_0,
  input         io_in_1,
  input         io_in_2,
  input         io_in_3,
  output        io_outR,
  output        io_outT,
  input         io_gndOuts,
  input         io_clkEnb
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] lut_in; // @[CLBlut4N10Clb.scala 73:27]
  wire [3:0] lut_sel; // @[CLBlut4N10Clb.scala 73:27]
  wire  lut_o; // @[CLBlut4N10Clb.scala 73:27]
  wire [1:0] lut_io_sel_lo = {io_in_1,io_in_0}; // @[CLBlut4N10Clb.scala 75:23]
  wire [1:0] lut_io_sel_hi = {io_in_3,io_in_2}; // @[CLBlut4N10Clb.scala 75:23]
  wire  _bleFF_T = ~io_clkEnb; // @[CLBlut4N10Clb.scala 77:48]
  reg  bleFF; // @[Reg.scala 28:20]
  wire  _io_outR_T_1 = io_config[16] ? lut_o : bleFF; // @[CLBlut4N10Clb.scala 80:17]
  wire  _io_outR_T_2 = ~io_gndOuts; // @[CLBlut4N10Clb.scala 80:52]
  wire  _io_outT_T_1 = io_config[17] ? lut_o : bleFF; // @[CLBlut4N10Clb.scala 81:17]
  Mux16C lut ( // @[CLBlut4N10Clb.scala 73:27]
    .in(lut_in),
    .sel(lut_sel),
    .o(lut_o)
  );
  assign io_outR = _io_outR_T_1 & ~io_gndOuts; // @[CLBlut4N10Clb.scala 80:50]
  assign io_outT = _io_outT_T_1 & _io_outR_T_2; // @[CLBlut4N10Clb.scala 81:50]
  assign lut_in = io_config[15:0]; // @[CLBlut4N10Clb.scala 74:25]
  assign lut_sel = {lut_io_sel_hi,lut_io_sel_lo}; // @[CLBlut4N10Clb.scala 75:23]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      bleFF <= 1'h0; // @[Reg.scala 28:20]
    end else if (_bleFF_T) begin // @[Reg.scala 29:18]
      bleFF <= lut_o; // @[Reg.scala 29:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bleFF = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLBlut4N10Alu(
  input          IPIN_0,
  input          IPIN_1,
  input          IPIN_2,
  input          IPIN_3,
  input          IPIN_4,
  input          IPIN_5,
  input          IPIN_6,
  input          IPIN_7,
  input          IPIN_8,
  input          IPIN_9,
  input          IPIN_10,
  input          IPIN_11,
  input          IPIN_12,
  input          IPIN_13,
  input          IPIN_14,
  input          IPIN_15,
  input          IPIN_16,
  input          IPIN_17,
  input          IPIN_18,
  input          IPIN_19,
  input          IPIN_20,
  input          IPIN_21,
  input          IPIN_22,
  input          IPIN_23,
  input          IPIN_24,
  input          IPIN_25,
  input          IPIN_26,
  input          IPIN_27,
  input          IPIN_28,
  input          IPIN_29,
  input          IPIN_30,
  input          IPIN_31,
  input          IPIN_32,
  input          IPIN_33,
  input          IPIN_34,
  input          IPIN_35,
  input          IPIN_36,
  input          IPIN_37,
  input          IPIN_38,
  input          IPIN_39,
  input          IPIN_40,
  input          IPIN_41,
  input          IPIN_42,
  input          IPIN_43,
  input          IPIN_44,
  input          IPIN_45,
  input          IPIN_46,
  input          IPIN_47,
  input          IPIN_48,
  input          IPIN_49,
  input          IPIN_50,
  input          IPIN_51,
  input          IPIN_52,
  input          IPIN_53,
  input          IPIN_54,
  input          IPIN_55,
  input          IPIN_56,
  input          IPIN_57,
  input          IPIN_58,
  input          IPIN_59,
  input          IPIN_60,
  input          IPIN_61,
  input          IPIN_62,
  input          IPIN_63,
  input          IPIN_64,
  input          IPIN_65,
  input          IPIN_66,
  input          IPIN_67,
  input          IPIN_68,
  input          IPIN_69,
  input          IPIN_70,
  input          IPIN_71,
  output         OPIN_73,
  output         OPIN_74,
  output         OPIN_75,
  output         OPIN_76,
  output         OPIN_77,
  output         OPIN_78,
  output         OPIN_79,
  output         OPIN_80,
  output         OPIN_81,
  output         OPIN_82,
  output         OPIN_83,
  output         OPIN_84,
  output         OPIN_85,
  output         OPIN_86,
  output         OPIN_87,
  output         OPIN_88,
  output         OPIN_89,
  output         OPIN_90,
  output         OPIN_91,
  output         OPIN_92,
  output         OPIN_93,
  output         OPIN_94,
  output         OPIN_95,
  output         OPIN_96,
  output         OPIN_97,
  output         OPIN_98,
  output         OPIN_99,
  output         OPIN_100,
  output         OPIN_101,
  output         OPIN_102,
  output         OPIN_103,
  output         OPIN_104,
  output         OPIN_105,
  output         OPIN_106,
  output         OPIN_107,
  output         OPIN_108,
  output         OPIN_109,
  output         OPIN_110,
  output         OPIN_111,
  output         OPIN_112,
  output         OPIN_113,
  output         OPIN_114,
  output         OPIN_115,
  output         OPIN_116,
  output         OPIN_117,
  output         OPIN_118,
  output         OPIN_119,
  output         OPIN_120,
  input          clock,
  input          reset,
  input  [193:0] configBits,
  input          gndLBouts
);
  wire  alu_clock; // @[CLBlut4N10Alu.scala 45:53]
  wire  alu_reset; // @[CLBlut4N10Alu.scala 45:53]
  wire [15:0] alu_io_i0; // @[CLBlut4N10Alu.scala 45:53]
  wire [15:0] alu_io_i1; // @[CLBlut4N10Alu.scala 45:53]
  wire [31:0] alu_io_ib32; // @[CLBlut4N10Alu.scala 45:53]
  wire [7:0] alu_io_ctrl; // @[CLBlut4N10Alu.scala 45:53]
  wire [15:0] alu_io_q; // @[CLBlut4N10Alu.scala 45:53]
  wire [31:0] alu_io_ob32; // @[CLBlut4N10Alu.scala 45:53]
  wire [31:0] alu_io_config; // @[CLBlut4N10Alu.scala 45:53]
  wire  alu_io_gndOuts; // @[CLBlut4N10Alu.scala 45:53]
  wire  alu_io_clkEnb; // @[CLBlut4N10Alu.scala 45:53]
  wire  BLE_0_clock; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_0_reset; // @[CLBlut4N10Alu.scala 64:48]
  wire [19:0] BLE_0_io_config; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_0_io_in_0; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_0_io_in_1; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_0_io_in_2; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_0_io_in_3; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_0_io_outR; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_0_io_outT; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_0_io_gndOuts; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_0_io_clkEnb; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_1_clock; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_1_reset; // @[CLBlut4N10Alu.scala 64:48]
  wire [19:0] BLE_1_io_config; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_1_io_in_0; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_1_io_in_1; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_1_io_in_2; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_1_io_in_3; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_1_io_outR; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_1_io_outT; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_1_io_gndOuts; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_1_io_clkEnb; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_2_clock; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_2_reset; // @[CLBlut4N10Alu.scala 64:48]
  wire [19:0] BLE_2_io_config; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_2_io_in_0; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_2_io_in_1; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_2_io_in_2; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_2_io_in_3; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_2_io_outR; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_2_io_outT; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_2_io_gndOuts; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_2_io_clkEnb; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_3_clock; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_3_reset; // @[CLBlut4N10Alu.scala 64:48]
  wire [19:0] BLE_3_io_config; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_3_io_in_0; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_3_io_in_1; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_3_io_in_2; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_3_io_in_3; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_3_io_outR; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_3_io_outT; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_3_io_gndOuts; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_3_io_clkEnb; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_4_clock; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_4_reset; // @[CLBlut4N10Alu.scala 64:48]
  wire [19:0] BLE_4_io_config; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_4_io_in_0; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_4_io_in_1; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_4_io_in_2; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_4_io_in_3; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_4_io_outR; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_4_io_outT; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_4_io_gndOuts; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_4_io_clkEnb; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_5_clock; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_5_reset; // @[CLBlut4N10Alu.scala 64:48]
  wire [19:0] BLE_5_io_config; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_5_io_in_0; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_5_io_in_1; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_5_io_in_2; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_5_io_in_3; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_5_io_outR; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_5_io_outT; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_5_io_gndOuts; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_5_io_clkEnb; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_6_clock; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_6_reset; // @[CLBlut4N10Alu.scala 64:48]
  wire [19:0] BLE_6_io_config; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_6_io_in_0; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_6_io_in_1; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_6_io_in_2; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_6_io_in_3; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_6_io_outR; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_6_io_outT; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_6_io_gndOuts; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_6_io_clkEnb; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_7_clock; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_7_reset; // @[CLBlut4N10Alu.scala 64:48]
  wire [19:0] BLE_7_io_config; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_7_io_in_0; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_7_io_in_1; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_7_io_in_2; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_7_io_in_3; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_7_io_outR; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_7_io_outT; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_7_io_gndOuts; // @[CLBlut4N10Alu.scala 64:48]
  wire  BLE_7_io_clkEnb; // @[CLBlut4N10Alu.scala 64:48]
  wire [7:0] I_0 = {IPIN_7,IPIN_6,IPIN_5,IPIN_4,IPIN_3,IPIN_2,IPIN_1,IPIN_0}; // @[CLBlut4N10Alu.scala 35:92]
  wire [7:0] I_1 = {IPIN_15,IPIN_14,IPIN_13,IPIN_12,IPIN_11,IPIN_10,IPIN_9,IPIN_8}; // @[CLBlut4N10Alu.scala 35:92]
  wire [7:0] I_2 = {IPIN_23,IPIN_22,IPIN_21,IPIN_20,IPIN_19,IPIN_18,IPIN_17,IPIN_16}; // @[CLBlut4N10Alu.scala 35:92]
  wire [7:0] I_3 = {IPIN_31,IPIN_30,IPIN_29,IPIN_28,IPIN_27,IPIN_26,IPIN_25,IPIN_24}; // @[CLBlut4N10Alu.scala 35:92]
  wire  OAlu_0 = alu_io_q[0]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_0 = BLE_0_io_outR; // @[CLBlut4N10Alu.scala 38:18 68:15]
  wire  OAlu_1 = alu_io_q[1]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_1 = BLE_1_io_outR; // @[CLBlut4N10Alu.scala 38:18 68:15]
  wire  OAlu_2 = alu_io_q[2]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_2 = BLE_2_io_outR; // @[CLBlut4N10Alu.scala 38:18 68:15]
  wire  OAlu_3 = alu_io_q[3]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_3 = BLE_3_io_outR; // @[CLBlut4N10Alu.scala 38:18 68:15]
  wire  OAlu_4 = alu_io_q[4]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_4 = BLE_4_io_outR; // @[CLBlut4N10Alu.scala 38:18 68:15]
  wire  OAlu_5 = alu_io_q[5]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_5 = BLE_5_io_outR; // @[CLBlut4N10Alu.scala 38:18 68:15]
  wire  OAlu_6 = alu_io_q[6]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_6 = BLE_6_io_outR; // @[CLBlut4N10Alu.scala 38:18 68:15]
  wire  OAlu_7 = alu_io_q[7]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_7 = BLE_7_io_outR; // @[CLBlut4N10Alu.scala 38:18 68:15]
  wire  OAlu_8 = alu_io_q[8]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_8 = BLE_0_io_outT; // @[CLBlut4N10Alu.scala 38:18 69:17]
  wire  OAlu_9 = alu_io_q[9]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_9 = BLE_1_io_outT; // @[CLBlut4N10Alu.scala 38:18 69:17]
  wire  OAlu_10 = alu_io_q[10]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_10 = BLE_2_io_outT; // @[CLBlut4N10Alu.scala 38:18 69:17]
  wire  OAlu_11 = alu_io_q[11]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_11 = BLE_3_io_outT; // @[CLBlut4N10Alu.scala 38:18 69:17]
  wire  OAlu_12 = alu_io_q[12]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_12 = BLE_4_io_outT; // @[CLBlut4N10Alu.scala 38:18 69:17]
  wire  OAlu_13 = alu_io_q[13]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_13 = BLE_5_io_outT; // @[CLBlut4N10Alu.scala 38:18 69:17]
  wire  OAlu_14 = alu_io_q[14]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_14 = BLE_6_io_outT; // @[CLBlut4N10Alu.scala 38:18 69:17]
  wire  OAlu_15 = alu_io_q[15]; // @[CLBlut4N10Alu.scala 50:50]
  wire  OClb_15 = BLE_7_io_outT; // @[CLBlut4N10Alu.scala 38:18 69:17]
  wire  OAlu_16 = alu_io_ob32[0]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_17 = alu_io_ob32[1]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_18 = alu_io_ob32[2]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_19 = alu_io_ob32[3]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_20 = alu_io_ob32[4]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_21 = alu_io_ob32[5]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_22 = alu_io_ob32[6]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_23 = alu_io_ob32[7]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_24 = alu_io_ob32[8]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_25 = alu_io_ob32[9]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_26 = alu_io_ob32[10]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_27 = alu_io_ob32[11]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_28 = alu_io_ob32[12]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_29 = alu_io_ob32[13]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_30 = alu_io_ob32[14]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_31 = alu_io_ob32[15]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_32 = alu_io_ob32[16]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_33 = alu_io_ob32[17]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_34 = alu_io_ob32[18]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_35 = alu_io_ob32[19]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_36 = alu_io_ob32[20]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_37 = alu_io_ob32[21]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_38 = alu_io_ob32[22]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_39 = alu_io_ob32[23]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_40 = alu_io_ob32[24]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_41 = alu_io_ob32[25]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_42 = alu_io_ob32[26]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_43 = alu_io_ob32[27]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_44 = alu_io_ob32[28]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_45 = alu_io_ob32[29]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_46 = alu_io_ob32[30]; // @[CLBlut4N10Alu.scala 51:54]
  wire  OAlu_47 = alu_io_ob32[31]; // @[CLBlut4N10Alu.scala 51:54]
  wire [8:0] IPINsasUint_lo_lo_lo = {IPIN_8,IPIN_7,IPIN_6,IPIN_5,IPIN_4,IPIN_3,IPIN_2,IPIN_1,IPIN_0}; // @[CLBlut4N10Alu.scala 44:50]
  wire [17:0] IPINsasUint_lo_lo = {IPIN_17,IPIN_16,IPIN_15,IPIN_14,IPIN_13,IPIN_12,IPIN_11,IPIN_10,IPIN_9,
    IPINsasUint_lo_lo_lo}; // @[CLBlut4N10Alu.scala 44:50]
  wire [8:0] IPINsasUint_lo_hi_lo = {IPIN_26,IPIN_25,IPIN_24,IPIN_23,IPIN_22,IPIN_21,IPIN_20,IPIN_19,IPIN_18}; // @[CLBlut4N10Alu.scala 44:50]
  wire [17:0] IPINsasUint_lo_hi = {IPIN_35,IPIN_34,IPIN_33,IPIN_32,IPIN_31,IPIN_30,IPIN_29,IPIN_28,IPIN_27,
    IPINsasUint_lo_hi_lo}; // @[CLBlut4N10Alu.scala 44:50]
  wire [8:0] IPINsasUint_hi_lo_lo = {IPIN_44,IPIN_43,IPIN_42,IPIN_41,IPIN_40,IPIN_39,IPIN_38,IPIN_37,IPIN_36}; // @[CLBlut4N10Alu.scala 44:50]
  wire [17:0] IPINsasUint_hi_lo = {IPIN_53,IPIN_52,IPIN_51,IPIN_50,IPIN_49,IPIN_48,IPIN_47,IPIN_46,IPIN_45,
    IPINsasUint_hi_lo_lo}; // @[CLBlut4N10Alu.scala 44:50]
  wire [8:0] IPINsasUint_hi_hi_lo = {IPIN_62,IPIN_61,IPIN_60,IPIN_59,IPIN_58,IPIN_57,IPIN_56,IPIN_55,IPIN_54}; // @[CLBlut4N10Alu.scala 44:50]
  wire [17:0] IPINsasUint_hi_hi = {IPIN_71,IPIN_70,IPIN_69,IPIN_68,IPIN_67,IPIN_66,IPIN_65,IPIN_64,IPIN_63,
    IPINsasUint_hi_hi_lo}; // @[CLBlut4N10Alu.scala 44:50]
  wire [71:0] IPINsasUint = {IPINsasUint_hi_hi,IPINsasUint_hi_lo,IPINsasUint_lo_hi,IPINsasUint_lo_lo}; // @[CLBlut4N10Alu.scala 44:50]
  Alu alu ( // @[CLBlut4N10Alu.scala 45:53]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_i0(alu_io_i0),
    .io_i1(alu_io_i1),
    .io_ib32(alu_io_ib32),
    .io_ctrl(alu_io_ctrl),
    .io_q(alu_io_q),
    .io_ob32(alu_io_ob32),
    .io_config(alu_io_config),
    .io_gndOuts(alu_io_gndOuts),
    .io_clkEnb(alu_io_clkEnb)
  );
  Ble4 BLE_0 ( // @[CLBlut4N10Alu.scala 64:48]
    .clock(BLE_0_clock),
    .reset(BLE_0_reset),
    .io_config(BLE_0_io_config),
    .io_in_0(BLE_0_io_in_0),
    .io_in_1(BLE_0_io_in_1),
    .io_in_2(BLE_0_io_in_2),
    .io_in_3(BLE_0_io_in_3),
    .io_outR(BLE_0_io_outR),
    .io_outT(BLE_0_io_outT),
    .io_gndOuts(BLE_0_io_gndOuts),
    .io_clkEnb(BLE_0_io_clkEnb)
  );
  Ble4 BLE_1 ( // @[CLBlut4N10Alu.scala 64:48]
    .clock(BLE_1_clock),
    .reset(BLE_1_reset),
    .io_config(BLE_1_io_config),
    .io_in_0(BLE_1_io_in_0),
    .io_in_1(BLE_1_io_in_1),
    .io_in_2(BLE_1_io_in_2),
    .io_in_3(BLE_1_io_in_3),
    .io_outR(BLE_1_io_outR),
    .io_outT(BLE_1_io_outT),
    .io_gndOuts(BLE_1_io_gndOuts),
    .io_clkEnb(BLE_1_io_clkEnb)
  );
  Ble4 BLE_2 ( // @[CLBlut4N10Alu.scala 64:48]
    .clock(BLE_2_clock),
    .reset(BLE_2_reset),
    .io_config(BLE_2_io_config),
    .io_in_0(BLE_2_io_in_0),
    .io_in_1(BLE_2_io_in_1),
    .io_in_2(BLE_2_io_in_2),
    .io_in_3(BLE_2_io_in_3),
    .io_outR(BLE_2_io_outR),
    .io_outT(BLE_2_io_outT),
    .io_gndOuts(BLE_2_io_gndOuts),
    .io_clkEnb(BLE_2_io_clkEnb)
  );
  Ble4 BLE_3 ( // @[CLBlut4N10Alu.scala 64:48]
    .clock(BLE_3_clock),
    .reset(BLE_3_reset),
    .io_config(BLE_3_io_config),
    .io_in_0(BLE_3_io_in_0),
    .io_in_1(BLE_3_io_in_1),
    .io_in_2(BLE_3_io_in_2),
    .io_in_3(BLE_3_io_in_3),
    .io_outR(BLE_3_io_outR),
    .io_outT(BLE_3_io_outT),
    .io_gndOuts(BLE_3_io_gndOuts),
    .io_clkEnb(BLE_3_io_clkEnb)
  );
  Ble4 BLE_4 ( // @[CLBlut4N10Alu.scala 64:48]
    .clock(BLE_4_clock),
    .reset(BLE_4_reset),
    .io_config(BLE_4_io_config),
    .io_in_0(BLE_4_io_in_0),
    .io_in_1(BLE_4_io_in_1),
    .io_in_2(BLE_4_io_in_2),
    .io_in_3(BLE_4_io_in_3),
    .io_outR(BLE_4_io_outR),
    .io_outT(BLE_4_io_outT),
    .io_gndOuts(BLE_4_io_gndOuts),
    .io_clkEnb(BLE_4_io_clkEnb)
  );
  Ble4 BLE_5 ( // @[CLBlut4N10Alu.scala 64:48]
    .clock(BLE_5_clock),
    .reset(BLE_5_reset),
    .io_config(BLE_5_io_config),
    .io_in_0(BLE_5_io_in_0),
    .io_in_1(BLE_5_io_in_1),
    .io_in_2(BLE_5_io_in_2),
    .io_in_3(BLE_5_io_in_3),
    .io_outR(BLE_5_io_outR),
    .io_outT(BLE_5_io_outT),
    .io_gndOuts(BLE_5_io_gndOuts),
    .io_clkEnb(BLE_5_io_clkEnb)
  );
  Ble4 BLE_6 ( // @[CLBlut4N10Alu.scala 64:48]
    .clock(BLE_6_clock),
    .reset(BLE_6_reset),
    .io_config(BLE_6_io_config),
    .io_in_0(BLE_6_io_in_0),
    .io_in_1(BLE_6_io_in_1),
    .io_in_2(BLE_6_io_in_2),
    .io_in_3(BLE_6_io_in_3),
    .io_outR(BLE_6_io_outR),
    .io_outT(BLE_6_io_outT),
    .io_gndOuts(BLE_6_io_gndOuts),
    .io_clkEnb(BLE_6_io_clkEnb)
  );
  Ble4 BLE_7 ( // @[CLBlut4N10Alu.scala 64:48]
    .clock(BLE_7_clock),
    .reset(BLE_7_reset),
    .io_config(BLE_7_io_config),
    .io_in_0(BLE_7_io_in_0),
    .io_in_1(BLE_7_io_in_1),
    .io_in_2(BLE_7_io_in_2),
    .io_in_3(BLE_7_io_in_3),
    .io_outR(BLE_7_io_outR),
    .io_outT(BLE_7_io_outT),
    .io_gndOuts(BLE_7_io_gndOuts),
    .io_clkEnb(BLE_7_io_clkEnb)
  );
  assign OPIN_73 = configBits[192] ? OAlu_0 & ~gndLBouts : OClb_0; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_74 = configBits[192] ? OAlu_1 & ~gndLBouts : OClb_1; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_75 = configBits[192] ? OAlu_2 & ~gndLBouts : OClb_2; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_76 = configBits[192] ? OAlu_3 & ~gndLBouts : OClb_3; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_77 = configBits[192] ? OAlu_4 & ~gndLBouts : OClb_4; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_78 = configBits[192] ? OAlu_5 & ~gndLBouts : OClb_5; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_79 = configBits[192] ? OAlu_6 & ~gndLBouts : OClb_6; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_80 = configBits[192] ? OAlu_7 & ~gndLBouts : OClb_7; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_81 = configBits[192] ? OAlu_8 & ~gndLBouts : OClb_8; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_82 = configBits[192] ? OAlu_9 & ~gndLBouts : OClb_9; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_83 = configBits[192] ? OAlu_10 & ~gndLBouts : OClb_10; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_84 = configBits[192] ? OAlu_11 & ~gndLBouts : OClb_11; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_85 = configBits[192] ? OAlu_12 & ~gndLBouts : OClb_12; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_86 = configBits[192] ? OAlu_13 & ~gndLBouts : OClb_13; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_87 = configBits[192] ? OAlu_14 & ~gndLBouts : OClb_14; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_88 = configBits[192] ? OAlu_15 & ~gndLBouts : OClb_15; // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_89 = configBits[192] & (OAlu_16 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_90 = configBits[192] & (OAlu_17 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_91 = configBits[192] & (OAlu_18 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_92 = configBits[192] & (OAlu_19 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_93 = configBits[192] & (OAlu_20 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_94 = configBits[192] & (OAlu_21 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_95 = configBits[192] & (OAlu_22 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_96 = configBits[192] & (OAlu_23 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_97 = configBits[192] & (OAlu_24 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_98 = configBits[192] & (OAlu_25 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_99 = configBits[192] & (OAlu_26 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_100 = configBits[192] & (OAlu_27 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_101 = configBits[192] & (OAlu_28 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_102 = configBits[192] & (OAlu_29 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_103 = configBits[192] & (OAlu_30 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_104 = configBits[192] & (OAlu_31 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_105 = configBits[192] & (OAlu_32 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_106 = configBits[192] & (OAlu_33 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_107 = configBits[192] & (OAlu_34 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_108 = configBits[192] & (OAlu_35 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_109 = configBits[192] & (OAlu_36 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_110 = configBits[192] & (OAlu_37 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_111 = configBits[192] & (OAlu_38 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_112 = configBits[192] & (OAlu_39 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_113 = configBits[192] & (OAlu_40 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_114 = configBits[192] & (OAlu_41 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_115 = configBits[192] & (OAlu_42 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_116 = configBits[192] & (OAlu_43 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_117 = configBits[192] & (OAlu_44 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_118 = configBits[192] & (OAlu_45 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_119 = configBits[192] & (OAlu_46 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign OPIN_120 = configBits[192] & (OAlu_47 & ~gndLBouts); // @[CLBlut4N10Alu.scala 40:15]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_i0 = IPINsasUint[15:0]; // @[CLBlut4N10Alu.scala 46:27]
  assign alu_io_i1 = IPINsasUint[31:16]; // @[CLBlut4N10Alu.scala 47:27]
  assign alu_io_ib32 = IPINsasUint[71:40]; // @[CLBlut4N10Alu.scala 49:29]
  assign alu_io_ctrl = IPINsasUint[39:32]; // @[CLBlut4N10Alu.scala 48:29]
  assign alu_io_config = configBits[33:2]; // @[CLBlut4N10Alu.scala 54:30]
  assign alu_io_gndOuts = gndLBouts; // @[CLBlut4N10Alu.scala 53:18]
  assign alu_io_clkEnb = configBits[193]; // @[CLBlut4N10Alu.scala 52:30]
  assign BLE_0_clock = clock;
  assign BLE_0_reset = reset;
  assign BLE_0_io_config = configBits[19:0]; // @[CLBlut4N10Alu.scala 66:38]
  assign BLE_0_io_in_0 = I_0[0]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_0_io_in_1 = I_1[0]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_0_io_in_2 = I_2[0]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_0_io_in_3 = I_3[0]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_0_io_gndOuts = gndLBouts; // @[CLBlut4N10Alu.scala 70:26]
  assign BLE_0_io_clkEnb = configBits[193]; // @[CLBlut4N10Alu.scala 71:38]
  assign BLE_1_clock = clock;
  assign BLE_1_reset = reset;
  assign BLE_1_io_config = configBits[39:20]; // @[CLBlut4N10Alu.scala 66:38]
  assign BLE_1_io_in_0 = I_0[1]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_1_io_in_1 = I_1[1]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_1_io_in_2 = I_2[1]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_1_io_in_3 = I_3[1]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_1_io_gndOuts = gndLBouts; // @[CLBlut4N10Alu.scala 70:26]
  assign BLE_1_io_clkEnb = configBits[193]; // @[CLBlut4N10Alu.scala 71:38]
  assign BLE_2_clock = clock;
  assign BLE_2_reset = reset;
  assign BLE_2_io_config = configBits[59:40]; // @[CLBlut4N10Alu.scala 66:38]
  assign BLE_2_io_in_0 = I_0[2]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_2_io_in_1 = I_1[2]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_2_io_in_2 = I_2[2]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_2_io_in_3 = I_3[2]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_2_io_gndOuts = gndLBouts; // @[CLBlut4N10Alu.scala 70:26]
  assign BLE_2_io_clkEnb = configBits[193]; // @[CLBlut4N10Alu.scala 71:38]
  assign BLE_3_clock = clock;
  assign BLE_3_reset = reset;
  assign BLE_3_io_config = configBits[79:60]; // @[CLBlut4N10Alu.scala 66:38]
  assign BLE_3_io_in_0 = I_0[3]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_3_io_in_1 = I_1[3]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_3_io_in_2 = I_2[3]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_3_io_in_3 = I_3[3]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_3_io_gndOuts = gndLBouts; // @[CLBlut4N10Alu.scala 70:26]
  assign BLE_3_io_clkEnb = configBits[193]; // @[CLBlut4N10Alu.scala 71:38]
  assign BLE_4_clock = clock;
  assign BLE_4_reset = reset;
  assign BLE_4_io_config = configBits[99:80]; // @[CLBlut4N10Alu.scala 66:38]
  assign BLE_4_io_in_0 = I_0[4]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_4_io_in_1 = I_1[4]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_4_io_in_2 = I_2[4]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_4_io_in_3 = I_3[4]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_4_io_gndOuts = gndLBouts; // @[CLBlut4N10Alu.scala 70:26]
  assign BLE_4_io_clkEnb = configBits[193]; // @[CLBlut4N10Alu.scala 71:38]
  assign BLE_5_clock = clock;
  assign BLE_5_reset = reset;
  assign BLE_5_io_config = configBits[119:100]; // @[CLBlut4N10Alu.scala 66:38]
  assign BLE_5_io_in_0 = I_0[5]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_5_io_in_1 = I_1[5]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_5_io_in_2 = I_2[5]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_5_io_in_3 = I_3[5]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_5_io_gndOuts = gndLBouts; // @[CLBlut4N10Alu.scala 70:26]
  assign BLE_5_io_clkEnb = configBits[193]; // @[CLBlut4N10Alu.scala 71:38]
  assign BLE_6_clock = clock;
  assign BLE_6_reset = reset;
  assign BLE_6_io_config = configBits[139:120]; // @[CLBlut4N10Alu.scala 66:38]
  assign BLE_6_io_in_0 = I_0[6]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_6_io_in_1 = I_1[6]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_6_io_in_2 = I_2[6]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_6_io_in_3 = I_3[6]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_6_io_gndOuts = gndLBouts; // @[CLBlut4N10Alu.scala 70:26]
  assign BLE_6_io_clkEnb = configBits[193]; // @[CLBlut4N10Alu.scala 71:38]
  assign BLE_7_clock = clock;
  assign BLE_7_reset = reset;
  assign BLE_7_io_config = configBits[159:140]; // @[CLBlut4N10Alu.scala 66:38]
  assign BLE_7_io_in_0 = I_0[7]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_7_io_in_1 = I_1[7]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_7_io_in_2 = I_2[7]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_7_io_in_3 = I_3[7]; // @[CLBlut4N10Alu.scala 67:62]
  assign BLE_7_io_gndOuts = gndLBouts; // @[CLBlut4N10Alu.scala 70:26]
  assign BLE_7_io_clkEnb = configBits[193]; // @[CLBlut4N10Alu.scala 71:38]
endmodule
module ScanConf_Tile_3_3_clbalutile(
  input          clock,
  output [511:0] ioBundle_confOut,
  input  [7:0]   ioBundle_scan_in,
  input          ioBundle_scan_en,
  output [7:0]   ioBundle_scan_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
`endif // RANDOMIZE_REG_INIT
  reg  confReg_0; // @[ScanConf.scala 32:20]
  reg  confReg_1; // @[ScanConf.scala 32:20]
  reg  confReg_2; // @[ScanConf.scala 32:20]
  reg  confReg_3; // @[ScanConf.scala 32:20]
  reg  confReg_4; // @[ScanConf.scala 32:20]
  reg  confReg_5; // @[ScanConf.scala 32:20]
  reg  confReg_6; // @[ScanConf.scala 32:20]
  reg  confReg_7; // @[ScanConf.scala 32:20]
  reg  confReg_8; // @[ScanConf.scala 32:20]
  reg  confReg_9; // @[ScanConf.scala 32:20]
  reg  confReg_10; // @[ScanConf.scala 32:20]
  reg  confReg_11; // @[ScanConf.scala 32:20]
  reg  confReg_12; // @[ScanConf.scala 32:20]
  reg  confReg_13; // @[ScanConf.scala 32:20]
  reg  confReg_14; // @[ScanConf.scala 32:20]
  reg  confReg_15; // @[ScanConf.scala 32:20]
  reg  confReg_16; // @[ScanConf.scala 32:20]
  reg  confReg_17; // @[ScanConf.scala 32:20]
  reg  confReg_18; // @[ScanConf.scala 32:20]
  reg  confReg_19; // @[ScanConf.scala 32:20]
  reg  confReg_20; // @[ScanConf.scala 32:20]
  reg  confReg_21; // @[ScanConf.scala 32:20]
  reg  confReg_22; // @[ScanConf.scala 32:20]
  reg  confReg_23; // @[ScanConf.scala 32:20]
  reg  confReg_24; // @[ScanConf.scala 32:20]
  reg  confReg_25; // @[ScanConf.scala 32:20]
  reg  confReg_26; // @[ScanConf.scala 32:20]
  reg  confReg_27; // @[ScanConf.scala 32:20]
  reg  confReg_28; // @[ScanConf.scala 32:20]
  reg  confReg_29; // @[ScanConf.scala 32:20]
  reg  confReg_30; // @[ScanConf.scala 32:20]
  reg  confReg_31; // @[ScanConf.scala 32:20]
  reg  confReg_32; // @[ScanConf.scala 32:20]
  reg  confReg_33; // @[ScanConf.scala 32:20]
  reg  confReg_34; // @[ScanConf.scala 32:20]
  reg  confReg_35; // @[ScanConf.scala 32:20]
  reg  confReg_36; // @[ScanConf.scala 32:20]
  reg  confReg_37; // @[ScanConf.scala 32:20]
  reg  confReg_38; // @[ScanConf.scala 32:20]
  reg  confReg_39; // @[ScanConf.scala 32:20]
  reg  confReg_40; // @[ScanConf.scala 32:20]
  reg  confReg_41; // @[ScanConf.scala 32:20]
  reg  confReg_42; // @[ScanConf.scala 32:20]
  reg  confReg_43; // @[ScanConf.scala 32:20]
  reg  confReg_44; // @[ScanConf.scala 32:20]
  reg  confReg_45; // @[ScanConf.scala 32:20]
  reg  confReg_46; // @[ScanConf.scala 32:20]
  reg  confReg_47; // @[ScanConf.scala 32:20]
  reg  confReg_48; // @[ScanConf.scala 32:20]
  reg  confReg_49; // @[ScanConf.scala 32:20]
  reg  confReg_50; // @[ScanConf.scala 32:20]
  reg  confReg_51; // @[ScanConf.scala 32:20]
  reg  confReg_52; // @[ScanConf.scala 32:20]
  reg  confReg_53; // @[ScanConf.scala 32:20]
  reg  confReg_54; // @[ScanConf.scala 32:20]
  reg  confReg_55; // @[ScanConf.scala 32:20]
  reg  confReg_56; // @[ScanConf.scala 32:20]
  reg  confReg_57; // @[ScanConf.scala 32:20]
  reg  confReg_58; // @[ScanConf.scala 32:20]
  reg  confReg_59; // @[ScanConf.scala 32:20]
  reg  confReg_60; // @[ScanConf.scala 32:20]
  reg  confReg_61; // @[ScanConf.scala 32:20]
  reg  confReg_62; // @[ScanConf.scala 32:20]
  reg  confReg_63; // @[ScanConf.scala 32:20]
  reg  confReg_64; // @[ScanConf.scala 32:20]
  reg  confReg_65; // @[ScanConf.scala 32:20]
  reg  confReg_66; // @[ScanConf.scala 32:20]
  reg  confReg_67; // @[ScanConf.scala 32:20]
  reg  confReg_68; // @[ScanConf.scala 32:20]
  reg  confReg_69; // @[ScanConf.scala 32:20]
  reg  confReg_70; // @[ScanConf.scala 32:20]
  reg  confReg_71; // @[ScanConf.scala 32:20]
  reg  confReg_72; // @[ScanConf.scala 32:20]
  reg  confReg_73; // @[ScanConf.scala 32:20]
  reg  confReg_74; // @[ScanConf.scala 32:20]
  reg  confReg_75; // @[ScanConf.scala 32:20]
  reg  confReg_76; // @[ScanConf.scala 32:20]
  reg  confReg_77; // @[ScanConf.scala 32:20]
  reg  confReg_78; // @[ScanConf.scala 32:20]
  reg  confReg_79; // @[ScanConf.scala 32:20]
  reg  confReg_80; // @[ScanConf.scala 32:20]
  reg  confReg_81; // @[ScanConf.scala 32:20]
  reg  confReg_82; // @[ScanConf.scala 32:20]
  reg  confReg_83; // @[ScanConf.scala 32:20]
  reg  confReg_84; // @[ScanConf.scala 32:20]
  reg  confReg_85; // @[ScanConf.scala 32:20]
  reg  confReg_86; // @[ScanConf.scala 32:20]
  reg  confReg_87; // @[ScanConf.scala 32:20]
  reg  confReg_88; // @[ScanConf.scala 32:20]
  reg  confReg_89; // @[ScanConf.scala 32:20]
  reg  confReg_90; // @[ScanConf.scala 32:20]
  reg  confReg_91; // @[ScanConf.scala 32:20]
  reg  confReg_92; // @[ScanConf.scala 32:20]
  reg  confReg_93; // @[ScanConf.scala 32:20]
  reg  confReg_94; // @[ScanConf.scala 32:20]
  reg  confReg_95; // @[ScanConf.scala 32:20]
  reg  confReg_96; // @[ScanConf.scala 32:20]
  reg  confReg_97; // @[ScanConf.scala 32:20]
  reg  confReg_98; // @[ScanConf.scala 32:20]
  reg  confReg_99; // @[ScanConf.scala 32:20]
  reg  confReg_100; // @[ScanConf.scala 32:20]
  reg  confReg_101; // @[ScanConf.scala 32:20]
  reg  confReg_102; // @[ScanConf.scala 32:20]
  reg  confReg_103; // @[ScanConf.scala 32:20]
  reg  confReg_104; // @[ScanConf.scala 32:20]
  reg  confReg_105; // @[ScanConf.scala 32:20]
  reg  confReg_106; // @[ScanConf.scala 32:20]
  reg  confReg_107; // @[ScanConf.scala 32:20]
  reg  confReg_108; // @[ScanConf.scala 32:20]
  reg  confReg_109; // @[ScanConf.scala 32:20]
  reg  confReg_110; // @[ScanConf.scala 32:20]
  reg  confReg_111; // @[ScanConf.scala 32:20]
  reg  confReg_112; // @[ScanConf.scala 32:20]
  reg  confReg_113; // @[ScanConf.scala 32:20]
  reg  confReg_114; // @[ScanConf.scala 32:20]
  reg  confReg_115; // @[ScanConf.scala 32:20]
  reg  confReg_116; // @[ScanConf.scala 32:20]
  reg  confReg_117; // @[ScanConf.scala 32:20]
  reg  confReg_118; // @[ScanConf.scala 32:20]
  reg  confReg_119; // @[ScanConf.scala 32:20]
  reg  confReg_120; // @[ScanConf.scala 32:20]
  reg  confReg_121; // @[ScanConf.scala 32:20]
  reg  confReg_122; // @[ScanConf.scala 32:20]
  reg  confReg_123; // @[ScanConf.scala 32:20]
  reg  confReg_124; // @[ScanConf.scala 32:20]
  reg  confReg_125; // @[ScanConf.scala 32:20]
  reg  confReg_126; // @[ScanConf.scala 32:20]
  reg  confReg_127; // @[ScanConf.scala 32:20]
  reg  confReg_128; // @[ScanConf.scala 32:20]
  reg  confReg_129; // @[ScanConf.scala 32:20]
  reg  confReg_130; // @[ScanConf.scala 32:20]
  reg  confReg_131; // @[ScanConf.scala 32:20]
  reg  confReg_132; // @[ScanConf.scala 32:20]
  reg  confReg_133; // @[ScanConf.scala 32:20]
  reg  confReg_134; // @[ScanConf.scala 32:20]
  reg  confReg_135; // @[ScanConf.scala 32:20]
  reg  confReg_136; // @[ScanConf.scala 32:20]
  reg  confReg_137; // @[ScanConf.scala 32:20]
  reg  confReg_138; // @[ScanConf.scala 32:20]
  reg  confReg_139; // @[ScanConf.scala 32:20]
  reg  confReg_140; // @[ScanConf.scala 32:20]
  reg  confReg_141; // @[ScanConf.scala 32:20]
  reg  confReg_142; // @[ScanConf.scala 32:20]
  reg  confReg_143; // @[ScanConf.scala 32:20]
  reg  confReg_144; // @[ScanConf.scala 32:20]
  reg  confReg_145; // @[ScanConf.scala 32:20]
  reg  confReg_146; // @[ScanConf.scala 32:20]
  reg  confReg_147; // @[ScanConf.scala 32:20]
  reg  confReg_148; // @[ScanConf.scala 32:20]
  reg  confReg_149; // @[ScanConf.scala 32:20]
  reg  confReg_150; // @[ScanConf.scala 32:20]
  reg  confReg_151; // @[ScanConf.scala 32:20]
  reg  confReg_152; // @[ScanConf.scala 32:20]
  reg  confReg_153; // @[ScanConf.scala 32:20]
  reg  confReg_154; // @[ScanConf.scala 32:20]
  reg  confReg_155; // @[ScanConf.scala 32:20]
  reg  confReg_156; // @[ScanConf.scala 32:20]
  reg  confReg_157; // @[ScanConf.scala 32:20]
  reg  confReg_158; // @[ScanConf.scala 32:20]
  reg  confReg_159; // @[ScanConf.scala 32:20]
  reg  confReg_160; // @[ScanConf.scala 32:20]
  reg  confReg_161; // @[ScanConf.scala 32:20]
  reg  confReg_162; // @[ScanConf.scala 32:20]
  reg  confReg_163; // @[ScanConf.scala 32:20]
  reg  confReg_164; // @[ScanConf.scala 32:20]
  reg  confReg_165; // @[ScanConf.scala 32:20]
  reg  confReg_166; // @[ScanConf.scala 32:20]
  reg  confReg_167; // @[ScanConf.scala 32:20]
  reg  confReg_168; // @[ScanConf.scala 32:20]
  reg  confReg_169; // @[ScanConf.scala 32:20]
  reg  confReg_170; // @[ScanConf.scala 32:20]
  reg  confReg_171; // @[ScanConf.scala 32:20]
  reg  confReg_172; // @[ScanConf.scala 32:20]
  reg  confReg_173; // @[ScanConf.scala 32:20]
  reg  confReg_174; // @[ScanConf.scala 32:20]
  reg  confReg_175; // @[ScanConf.scala 32:20]
  reg  confReg_176; // @[ScanConf.scala 32:20]
  reg  confReg_177; // @[ScanConf.scala 32:20]
  reg  confReg_178; // @[ScanConf.scala 32:20]
  reg  confReg_179; // @[ScanConf.scala 32:20]
  reg  confReg_180; // @[ScanConf.scala 32:20]
  reg  confReg_181; // @[ScanConf.scala 32:20]
  reg  confReg_182; // @[ScanConf.scala 32:20]
  reg  confReg_183; // @[ScanConf.scala 32:20]
  reg  confReg_184; // @[ScanConf.scala 32:20]
  reg  confReg_185; // @[ScanConf.scala 32:20]
  reg  confReg_186; // @[ScanConf.scala 32:20]
  reg  confReg_187; // @[ScanConf.scala 32:20]
  reg  confReg_188; // @[ScanConf.scala 32:20]
  reg  confReg_189; // @[ScanConf.scala 32:20]
  reg  confReg_190; // @[ScanConf.scala 32:20]
  reg  confReg_191; // @[ScanConf.scala 32:20]
  reg  confReg_192; // @[ScanConf.scala 32:20]
  reg  confReg_193; // @[ScanConf.scala 32:20]
  reg  confReg_194; // @[ScanConf.scala 32:20]
  reg  confReg_195; // @[ScanConf.scala 32:20]
  reg  confReg_196; // @[ScanConf.scala 32:20]
  reg  confReg_197; // @[ScanConf.scala 32:20]
  reg  confReg_198; // @[ScanConf.scala 32:20]
  reg  confReg_199; // @[ScanConf.scala 32:20]
  reg  confReg_200; // @[ScanConf.scala 32:20]
  reg  confReg_201; // @[ScanConf.scala 32:20]
  reg  confReg_202; // @[ScanConf.scala 32:20]
  reg  confReg_203; // @[ScanConf.scala 32:20]
  reg  confReg_204; // @[ScanConf.scala 32:20]
  reg  confReg_205; // @[ScanConf.scala 32:20]
  reg  confReg_206; // @[ScanConf.scala 32:20]
  reg  confReg_207; // @[ScanConf.scala 32:20]
  reg  confReg_208; // @[ScanConf.scala 32:20]
  reg  confReg_209; // @[ScanConf.scala 32:20]
  reg  confReg_210; // @[ScanConf.scala 32:20]
  reg  confReg_211; // @[ScanConf.scala 32:20]
  reg  confReg_212; // @[ScanConf.scala 32:20]
  reg  confReg_213; // @[ScanConf.scala 32:20]
  reg  confReg_214; // @[ScanConf.scala 32:20]
  reg  confReg_215; // @[ScanConf.scala 32:20]
  reg  confReg_216; // @[ScanConf.scala 32:20]
  reg  confReg_217; // @[ScanConf.scala 32:20]
  reg  confReg_218; // @[ScanConf.scala 32:20]
  reg  confReg_219; // @[ScanConf.scala 32:20]
  reg  confReg_220; // @[ScanConf.scala 32:20]
  reg  confReg_221; // @[ScanConf.scala 32:20]
  reg  confReg_222; // @[ScanConf.scala 32:20]
  reg  confReg_223; // @[ScanConf.scala 32:20]
  reg  confReg_224; // @[ScanConf.scala 32:20]
  reg  confReg_225; // @[ScanConf.scala 32:20]
  reg  confReg_226; // @[ScanConf.scala 32:20]
  reg  confReg_227; // @[ScanConf.scala 32:20]
  reg  confReg_228; // @[ScanConf.scala 32:20]
  reg  confReg_229; // @[ScanConf.scala 32:20]
  reg  confReg_230; // @[ScanConf.scala 32:20]
  reg  confReg_231; // @[ScanConf.scala 32:20]
  reg  confReg_232; // @[ScanConf.scala 32:20]
  reg  confReg_233; // @[ScanConf.scala 32:20]
  reg  confReg_234; // @[ScanConf.scala 32:20]
  reg  confReg_235; // @[ScanConf.scala 32:20]
  reg  confReg_236; // @[ScanConf.scala 32:20]
  reg  confReg_237; // @[ScanConf.scala 32:20]
  reg  confReg_238; // @[ScanConf.scala 32:20]
  reg  confReg_239; // @[ScanConf.scala 32:20]
  reg  confReg_240; // @[ScanConf.scala 32:20]
  reg  confReg_241; // @[ScanConf.scala 32:20]
  reg  confReg_242; // @[ScanConf.scala 32:20]
  reg  confReg_243; // @[ScanConf.scala 32:20]
  reg  confReg_244; // @[ScanConf.scala 32:20]
  reg  confReg_245; // @[ScanConf.scala 32:20]
  reg  confReg_246; // @[ScanConf.scala 32:20]
  reg  confReg_247; // @[ScanConf.scala 32:20]
  reg  confReg_248; // @[ScanConf.scala 32:20]
  reg  confReg_249; // @[ScanConf.scala 32:20]
  reg  confReg_250; // @[ScanConf.scala 32:20]
  reg  confReg_251; // @[ScanConf.scala 32:20]
  reg  confReg_252; // @[ScanConf.scala 32:20]
  reg  confReg_253; // @[ScanConf.scala 32:20]
  reg  confReg_254; // @[ScanConf.scala 32:20]
  reg  confReg_255; // @[ScanConf.scala 32:20]
  reg  confReg_256; // @[ScanConf.scala 32:20]
  reg  confReg_257; // @[ScanConf.scala 32:20]
  reg  confReg_258; // @[ScanConf.scala 32:20]
  reg  confReg_259; // @[ScanConf.scala 32:20]
  reg  confReg_260; // @[ScanConf.scala 32:20]
  reg  confReg_261; // @[ScanConf.scala 32:20]
  reg  confReg_262; // @[ScanConf.scala 32:20]
  reg  confReg_263; // @[ScanConf.scala 32:20]
  reg  confReg_264; // @[ScanConf.scala 32:20]
  reg  confReg_265; // @[ScanConf.scala 32:20]
  reg  confReg_266; // @[ScanConf.scala 32:20]
  reg  confReg_267; // @[ScanConf.scala 32:20]
  reg  confReg_268; // @[ScanConf.scala 32:20]
  reg  confReg_269; // @[ScanConf.scala 32:20]
  reg  confReg_270; // @[ScanConf.scala 32:20]
  reg  confReg_271; // @[ScanConf.scala 32:20]
  reg  confReg_272; // @[ScanConf.scala 32:20]
  reg  confReg_273; // @[ScanConf.scala 32:20]
  reg  confReg_274; // @[ScanConf.scala 32:20]
  reg  confReg_275; // @[ScanConf.scala 32:20]
  reg  confReg_276; // @[ScanConf.scala 32:20]
  reg  confReg_277; // @[ScanConf.scala 32:20]
  reg  confReg_278; // @[ScanConf.scala 32:20]
  reg  confReg_279; // @[ScanConf.scala 32:20]
  reg  confReg_280; // @[ScanConf.scala 32:20]
  reg  confReg_281; // @[ScanConf.scala 32:20]
  reg  confReg_282; // @[ScanConf.scala 32:20]
  reg  confReg_283; // @[ScanConf.scala 32:20]
  reg  confReg_284; // @[ScanConf.scala 32:20]
  reg  confReg_285; // @[ScanConf.scala 32:20]
  reg  confReg_286; // @[ScanConf.scala 32:20]
  reg  confReg_287; // @[ScanConf.scala 32:20]
  reg  confReg_288; // @[ScanConf.scala 32:20]
  reg  confReg_289; // @[ScanConf.scala 32:20]
  reg  confReg_290; // @[ScanConf.scala 32:20]
  reg  confReg_291; // @[ScanConf.scala 32:20]
  reg  confReg_292; // @[ScanConf.scala 32:20]
  reg  confReg_293; // @[ScanConf.scala 32:20]
  reg  confReg_294; // @[ScanConf.scala 32:20]
  reg  confReg_295; // @[ScanConf.scala 32:20]
  reg  confReg_296; // @[ScanConf.scala 32:20]
  reg  confReg_297; // @[ScanConf.scala 32:20]
  reg  confReg_298; // @[ScanConf.scala 32:20]
  reg  confReg_299; // @[ScanConf.scala 32:20]
  reg  confReg_300; // @[ScanConf.scala 32:20]
  reg  confReg_301; // @[ScanConf.scala 32:20]
  reg  confReg_302; // @[ScanConf.scala 32:20]
  reg  confReg_303; // @[ScanConf.scala 32:20]
  reg  confReg_304; // @[ScanConf.scala 32:20]
  reg  confReg_305; // @[ScanConf.scala 32:20]
  reg  confReg_306; // @[ScanConf.scala 32:20]
  reg  confReg_307; // @[ScanConf.scala 32:20]
  reg  confReg_308; // @[ScanConf.scala 32:20]
  reg  confReg_309; // @[ScanConf.scala 32:20]
  reg  confReg_310; // @[ScanConf.scala 32:20]
  reg  confReg_311; // @[ScanConf.scala 32:20]
  reg  confReg_312; // @[ScanConf.scala 32:20]
  reg  confReg_313; // @[ScanConf.scala 32:20]
  reg  confReg_314; // @[ScanConf.scala 32:20]
  reg  confReg_315; // @[ScanConf.scala 32:20]
  reg  confReg_316; // @[ScanConf.scala 32:20]
  reg  confReg_317; // @[ScanConf.scala 32:20]
  reg  confReg_318; // @[ScanConf.scala 32:20]
  reg  confReg_319; // @[ScanConf.scala 32:20]
  reg  confReg_320; // @[ScanConf.scala 32:20]
  reg  confReg_321; // @[ScanConf.scala 32:20]
  reg  confReg_322; // @[ScanConf.scala 32:20]
  reg  confReg_323; // @[ScanConf.scala 32:20]
  reg  confReg_324; // @[ScanConf.scala 32:20]
  reg  confReg_325; // @[ScanConf.scala 32:20]
  reg  confReg_326; // @[ScanConf.scala 32:20]
  reg  confReg_327; // @[ScanConf.scala 32:20]
  reg  confReg_328; // @[ScanConf.scala 32:20]
  reg  confReg_329; // @[ScanConf.scala 32:20]
  reg  confReg_330; // @[ScanConf.scala 32:20]
  reg  confReg_331; // @[ScanConf.scala 32:20]
  reg  confReg_332; // @[ScanConf.scala 32:20]
  reg  confReg_333; // @[ScanConf.scala 32:20]
  reg  confReg_334; // @[ScanConf.scala 32:20]
  reg  confReg_335; // @[ScanConf.scala 32:20]
  reg  confReg_336; // @[ScanConf.scala 32:20]
  reg  confReg_337; // @[ScanConf.scala 32:20]
  reg  confReg_338; // @[ScanConf.scala 32:20]
  reg  confReg_339; // @[ScanConf.scala 32:20]
  reg  confReg_340; // @[ScanConf.scala 32:20]
  reg  confReg_341; // @[ScanConf.scala 32:20]
  reg  confReg_342; // @[ScanConf.scala 32:20]
  reg  confReg_343; // @[ScanConf.scala 32:20]
  reg  confReg_344; // @[ScanConf.scala 32:20]
  reg  confReg_345; // @[ScanConf.scala 32:20]
  reg  confReg_346; // @[ScanConf.scala 32:20]
  reg  confReg_347; // @[ScanConf.scala 32:20]
  reg  confReg_348; // @[ScanConf.scala 32:20]
  reg  confReg_349; // @[ScanConf.scala 32:20]
  reg  confReg_350; // @[ScanConf.scala 32:20]
  reg  confReg_351; // @[ScanConf.scala 32:20]
  reg  confReg_352; // @[ScanConf.scala 32:20]
  reg  confReg_353; // @[ScanConf.scala 32:20]
  reg  confReg_354; // @[ScanConf.scala 32:20]
  reg  confReg_355; // @[ScanConf.scala 32:20]
  reg  confReg_356; // @[ScanConf.scala 32:20]
  reg  confReg_357; // @[ScanConf.scala 32:20]
  reg  confReg_358; // @[ScanConf.scala 32:20]
  reg  confReg_359; // @[ScanConf.scala 32:20]
  reg  confReg_360; // @[ScanConf.scala 32:20]
  reg  confReg_361; // @[ScanConf.scala 32:20]
  reg  confReg_362; // @[ScanConf.scala 32:20]
  reg  confReg_363; // @[ScanConf.scala 32:20]
  reg  confReg_364; // @[ScanConf.scala 32:20]
  reg  confReg_365; // @[ScanConf.scala 32:20]
  reg  confReg_366; // @[ScanConf.scala 32:20]
  reg  confReg_367; // @[ScanConf.scala 32:20]
  reg  confReg_368; // @[ScanConf.scala 32:20]
  reg  confReg_369; // @[ScanConf.scala 32:20]
  reg  confReg_370; // @[ScanConf.scala 32:20]
  reg  confReg_371; // @[ScanConf.scala 32:20]
  reg  confReg_372; // @[ScanConf.scala 32:20]
  reg  confReg_373; // @[ScanConf.scala 32:20]
  reg  confReg_374; // @[ScanConf.scala 32:20]
  reg  confReg_375; // @[ScanConf.scala 32:20]
  reg  confReg_376; // @[ScanConf.scala 32:20]
  reg  confReg_377; // @[ScanConf.scala 32:20]
  reg  confReg_378; // @[ScanConf.scala 32:20]
  reg  confReg_379; // @[ScanConf.scala 32:20]
  reg  confReg_380; // @[ScanConf.scala 32:20]
  reg  confReg_381; // @[ScanConf.scala 32:20]
  reg  confReg_382; // @[ScanConf.scala 32:20]
  reg  confReg_383; // @[ScanConf.scala 32:20]
  reg  confReg_384; // @[ScanConf.scala 32:20]
  reg  confReg_385; // @[ScanConf.scala 32:20]
  reg  confReg_386; // @[ScanConf.scala 32:20]
  reg  confReg_387; // @[ScanConf.scala 32:20]
  reg  confReg_388; // @[ScanConf.scala 32:20]
  reg  confReg_389; // @[ScanConf.scala 32:20]
  reg  confReg_390; // @[ScanConf.scala 32:20]
  reg  confReg_391; // @[ScanConf.scala 32:20]
  reg  confReg_392; // @[ScanConf.scala 32:20]
  reg  confReg_393; // @[ScanConf.scala 32:20]
  reg  confReg_394; // @[ScanConf.scala 32:20]
  reg  confReg_395; // @[ScanConf.scala 32:20]
  reg  confReg_396; // @[ScanConf.scala 32:20]
  reg  confReg_397; // @[ScanConf.scala 32:20]
  reg  confReg_398; // @[ScanConf.scala 32:20]
  reg  confReg_399; // @[ScanConf.scala 32:20]
  reg  confReg_400; // @[ScanConf.scala 32:20]
  reg  confReg_401; // @[ScanConf.scala 32:20]
  reg  confReg_402; // @[ScanConf.scala 32:20]
  reg  confReg_403; // @[ScanConf.scala 32:20]
  reg  confReg_404; // @[ScanConf.scala 32:20]
  reg  confReg_405; // @[ScanConf.scala 32:20]
  reg  confReg_406; // @[ScanConf.scala 32:20]
  reg  confReg_407; // @[ScanConf.scala 32:20]
  reg  confReg_408; // @[ScanConf.scala 32:20]
  reg  confReg_409; // @[ScanConf.scala 32:20]
  reg  confReg_410; // @[ScanConf.scala 32:20]
  reg  confReg_411; // @[ScanConf.scala 32:20]
  reg  confReg_412; // @[ScanConf.scala 32:20]
  reg  confReg_413; // @[ScanConf.scala 32:20]
  reg  confReg_414; // @[ScanConf.scala 32:20]
  reg  confReg_415; // @[ScanConf.scala 32:20]
  reg  confReg_416; // @[ScanConf.scala 32:20]
  reg  confReg_417; // @[ScanConf.scala 32:20]
  reg  confReg_418; // @[ScanConf.scala 32:20]
  reg  confReg_419; // @[ScanConf.scala 32:20]
  reg  confReg_420; // @[ScanConf.scala 32:20]
  reg  confReg_421; // @[ScanConf.scala 32:20]
  reg  confReg_422; // @[ScanConf.scala 32:20]
  reg  confReg_423; // @[ScanConf.scala 32:20]
  reg  confReg_424; // @[ScanConf.scala 32:20]
  reg  confReg_425; // @[ScanConf.scala 32:20]
  reg  confReg_426; // @[ScanConf.scala 32:20]
  reg  confReg_427; // @[ScanConf.scala 32:20]
  reg  confReg_428; // @[ScanConf.scala 32:20]
  reg  confReg_429; // @[ScanConf.scala 32:20]
  reg  confReg_430; // @[ScanConf.scala 32:20]
  reg  confReg_431; // @[ScanConf.scala 32:20]
  reg  confReg_432; // @[ScanConf.scala 32:20]
  reg  confReg_433; // @[ScanConf.scala 32:20]
  reg  confReg_434; // @[ScanConf.scala 32:20]
  reg  confReg_435; // @[ScanConf.scala 32:20]
  reg  confReg_436; // @[ScanConf.scala 32:20]
  reg  confReg_437; // @[ScanConf.scala 32:20]
  reg  confReg_438; // @[ScanConf.scala 32:20]
  reg  confReg_439; // @[ScanConf.scala 32:20]
  reg  confReg_440; // @[ScanConf.scala 32:20]
  reg  confReg_441; // @[ScanConf.scala 32:20]
  reg  confReg_442; // @[ScanConf.scala 32:20]
  reg  confReg_443; // @[ScanConf.scala 32:20]
  reg  confReg_444; // @[ScanConf.scala 32:20]
  reg  confReg_445; // @[ScanConf.scala 32:20]
  reg  confReg_446; // @[ScanConf.scala 32:20]
  reg  confReg_447; // @[ScanConf.scala 32:20]
  reg  confReg_448; // @[ScanConf.scala 32:20]
  reg  confReg_449; // @[ScanConf.scala 32:20]
  reg  confReg_450; // @[ScanConf.scala 32:20]
  reg  confReg_451; // @[ScanConf.scala 32:20]
  reg  confReg_452; // @[ScanConf.scala 32:20]
  reg  confReg_453; // @[ScanConf.scala 32:20]
  reg  confReg_454; // @[ScanConf.scala 32:20]
  reg  confReg_455; // @[ScanConf.scala 32:20]
  reg  confReg_456; // @[ScanConf.scala 32:20]
  reg  confReg_457; // @[ScanConf.scala 32:20]
  reg  confReg_458; // @[ScanConf.scala 32:20]
  reg  confReg_459; // @[ScanConf.scala 32:20]
  reg  confReg_460; // @[ScanConf.scala 32:20]
  reg  confReg_461; // @[ScanConf.scala 32:20]
  reg  confReg_462; // @[ScanConf.scala 32:20]
  reg  confReg_463; // @[ScanConf.scala 32:20]
  reg  confReg_464; // @[ScanConf.scala 32:20]
  reg  confReg_465; // @[ScanConf.scala 32:20]
  reg  confReg_466; // @[ScanConf.scala 32:20]
  reg  confReg_467; // @[ScanConf.scala 32:20]
  reg  confReg_468; // @[ScanConf.scala 32:20]
  reg  confReg_469; // @[ScanConf.scala 32:20]
  reg  confReg_470; // @[ScanConf.scala 32:20]
  reg  confReg_471; // @[ScanConf.scala 32:20]
  reg  confReg_472; // @[ScanConf.scala 32:20]
  reg  confReg_473; // @[ScanConf.scala 32:20]
  reg  confReg_474; // @[ScanConf.scala 32:20]
  reg  confReg_475; // @[ScanConf.scala 32:20]
  reg  confReg_476; // @[ScanConf.scala 32:20]
  reg  confReg_477; // @[ScanConf.scala 32:20]
  reg  confReg_478; // @[ScanConf.scala 32:20]
  reg  confReg_479; // @[ScanConf.scala 32:20]
  reg  confReg_480; // @[ScanConf.scala 32:20]
  reg  confReg_481; // @[ScanConf.scala 32:20]
  reg  confReg_482; // @[ScanConf.scala 32:20]
  reg  confReg_483; // @[ScanConf.scala 32:20]
  reg  confReg_484; // @[ScanConf.scala 32:20]
  reg  confReg_485; // @[ScanConf.scala 32:20]
  reg  confReg_486; // @[ScanConf.scala 32:20]
  reg  confReg_487; // @[ScanConf.scala 32:20]
  reg  confReg_488; // @[ScanConf.scala 32:20]
  reg  confReg_489; // @[ScanConf.scala 32:20]
  reg  confReg_490; // @[ScanConf.scala 32:20]
  reg  confReg_491; // @[ScanConf.scala 32:20]
  reg  confReg_492; // @[ScanConf.scala 32:20]
  reg  confReg_493; // @[ScanConf.scala 32:20]
  reg  confReg_494; // @[ScanConf.scala 32:20]
  reg  confReg_495; // @[ScanConf.scala 32:20]
  reg  confReg_496; // @[ScanConf.scala 32:20]
  reg  confReg_497; // @[ScanConf.scala 32:20]
  reg  confReg_498; // @[ScanConf.scala 32:20]
  reg  confReg_499; // @[ScanConf.scala 32:20]
  reg  confReg_500; // @[ScanConf.scala 32:20]
  reg  confReg_501; // @[ScanConf.scala 32:20]
  reg  confReg_502; // @[ScanConf.scala 32:20]
  reg  confReg_503; // @[ScanConf.scala 32:20]
  reg  confReg_504; // @[ScanConf.scala 32:20]
  reg  confReg_505; // @[ScanConf.scala 32:20]
  reg  confReg_506; // @[ScanConf.scala 32:20]
  reg  confReg_507; // @[ScanConf.scala 32:20]
  reg  confReg_508; // @[ScanConf.scala 32:20]
  reg  confReg_509; // @[ScanConf.scala 32:20]
  reg  confReg_510; // @[ScanConf.scala 32:20]
  reg  confReg_511; // @[ScanConf.scala 32:20]
  wire [3:0] io_scan_out_lo = {confReg_3,confReg_2,confReg_1,confReg_0}; // @[ScanConf.scala 46:47]
  wire [3:0] io_scan_out_hi = {confReg_7,confReg_6,confReg_5,confReg_4}; // @[ScanConf.scala 46:47]
  wire [7:0] io_scan_out = {confReg_7,confReg_6,confReg_5,confReg_4,confReg_3,confReg_2,confReg_1,confReg_0}; // @[ScanConf.scala 46:47]
  wire [15:0] io_confOut_lo_lo_lo_lo_lo = {confReg_15,confReg_14,confReg_13,confReg_12,confReg_11,confReg_10,confReg_9,
    confReg_8,io_scan_out}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_lo_lo_hi_lo = {confReg_23,confReg_22,confReg_21,confReg_20,confReg_19,confReg_18,
    confReg_17,confReg_16}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_lo_lo_lo = {confReg_31,confReg_30,confReg_29,confReg_28,confReg_27,confReg_26,confReg_25,
    confReg_24,io_confOut_lo_lo_lo_lo_hi_lo,io_confOut_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_lo_hi_lo_lo = {confReg_39,confReg_38,confReg_37,confReg_36,confReg_35,confReg_34,
    confReg_33,confReg_32}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_lo_lo_hi_lo = {confReg_47,confReg_46,confReg_45,confReg_44,confReg_43,confReg_42,confReg_41,
    confReg_40,io_confOut_lo_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_lo_hi_hi_lo = {confReg_55,confReg_54,confReg_53,confReg_52,confReg_51,confReg_50,
    confReg_49,confReg_48}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_lo_lo_hi = {confReg_63,confReg_62,confReg_61,confReg_60,confReg_59,confReg_58,confReg_57,
    confReg_56,io_confOut_lo_lo_lo_hi_hi_lo,io_confOut_lo_lo_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_hi_lo_lo_lo = {confReg_71,confReg_70,confReg_69,confReg_68,confReg_67,confReg_66,
    confReg_65,confReg_64}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_lo_hi_lo_lo = {confReg_79,confReg_78,confReg_77,confReg_76,confReg_75,confReg_74,confReg_73,
    confReg_72,io_confOut_lo_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_hi_lo_hi_lo = {confReg_87,confReg_86,confReg_85,confReg_84,confReg_83,confReg_82,
    confReg_81,confReg_80}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_lo_hi_lo = {confReg_95,confReg_94,confReg_93,confReg_92,confReg_91,confReg_90,confReg_89,
    confReg_88,io_confOut_lo_lo_hi_lo_hi_lo,io_confOut_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_hi_hi_lo_lo = {confReg_103,confReg_102,confReg_101,confReg_100,confReg_99,confReg_98,
    confReg_97,confReg_96}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_lo_hi_hi_lo = {confReg_111,confReg_110,confReg_109,confReg_108,confReg_107,confReg_106,
    confReg_105,confReg_104,io_confOut_lo_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_hi_hi_hi_lo = {confReg_119,confReg_118,confReg_117,confReg_116,confReg_115,confReg_114,
    confReg_113,confReg_112}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_lo_hi_hi = {confReg_127,confReg_126,confReg_125,confReg_124,confReg_123,confReg_122,
    confReg_121,confReg_120,io_confOut_lo_lo_hi_hi_hi_lo,io_confOut_lo_lo_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_lo_lo_lo_lo = {confReg_135,confReg_134,confReg_133,confReg_132,confReg_131,confReg_130,
    confReg_129,confReg_128}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_hi_lo_lo_lo = {confReg_143,confReg_142,confReg_141,confReg_140,confReg_139,confReg_138,
    confReg_137,confReg_136,io_confOut_lo_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_lo_lo_hi_lo = {confReg_151,confReg_150,confReg_149,confReg_148,confReg_147,confReg_146,
    confReg_145,confReg_144}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_hi_lo_lo = {confReg_159,confReg_158,confReg_157,confReg_156,confReg_155,confReg_154,
    confReg_153,confReg_152,io_confOut_lo_hi_lo_lo_hi_lo,io_confOut_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_lo_hi_lo_lo = {confReg_167,confReg_166,confReg_165,confReg_164,confReg_163,confReg_162,
    confReg_161,confReg_160}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_hi_lo_hi_lo = {confReg_175,confReg_174,confReg_173,confReg_172,confReg_171,confReg_170,
    confReg_169,confReg_168,io_confOut_lo_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_lo_hi_hi_lo = {confReg_183,confReg_182,confReg_181,confReg_180,confReg_179,confReg_178,
    confReg_177,confReg_176}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_hi_lo_hi = {confReg_191,confReg_190,confReg_189,confReg_188,confReg_187,confReg_186,
    confReg_185,confReg_184,io_confOut_lo_hi_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_hi_lo_lo_lo = {confReg_199,confReg_198,confReg_197,confReg_196,confReg_195,confReg_194,
    confReg_193,confReg_192}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_hi_hi_lo_lo = {confReg_207,confReg_206,confReg_205,confReg_204,confReg_203,confReg_202,
    confReg_201,confReg_200,io_confOut_lo_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_hi_lo_hi_lo = {confReg_215,confReg_214,confReg_213,confReg_212,confReg_211,confReg_210,
    confReg_209,confReg_208}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_hi_hi_lo = {confReg_223,confReg_222,confReg_221,confReg_220,confReg_219,confReg_218,
    confReg_217,confReg_216,io_confOut_lo_hi_hi_lo_hi_lo,io_confOut_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_hi_hi_lo_lo = {confReg_231,confReg_230,confReg_229,confReg_228,confReg_227,confReg_226,
    confReg_225,confReg_224}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_hi_hi_hi_lo = {confReg_239,confReg_238,confReg_237,confReg_236,confReg_235,confReg_234,
    confReg_233,confReg_232,io_confOut_lo_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_hi_hi_hi_lo = {confReg_247,confReg_246,confReg_245,confReg_244,confReg_243,confReg_242,
    confReg_241,confReg_240}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_hi_hi_hi = {confReg_255,confReg_254,confReg_253,confReg_252,confReg_251,confReg_250,
    confReg_249,confReg_248,io_confOut_lo_hi_hi_hi_hi_lo,io_confOut_lo_hi_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [255:0] io_confOut_lo = {io_confOut_lo_hi_hi_hi,io_confOut_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi,
    io_confOut_lo_hi_lo_lo,io_confOut_lo_lo_hi_hi,io_confOut_lo_lo_hi_lo,io_confOut_lo_lo_lo_hi,io_confOut_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_lo_lo_lo_lo = {confReg_263,confReg_262,confReg_261,confReg_260,confReg_259,confReg_258,
    confReg_257,confReg_256}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_lo_lo_lo_lo = {confReg_271,confReg_270,confReg_269,confReg_268,confReg_267,confReg_266,
    confReg_265,confReg_264,io_confOut_hi_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_lo_lo_hi_lo = {confReg_279,confReg_278,confReg_277,confReg_276,confReg_275,confReg_274,
    confReg_273,confReg_272}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_lo_lo_lo = {confReg_287,confReg_286,confReg_285,confReg_284,confReg_283,confReg_282,
    confReg_281,confReg_280,io_confOut_hi_lo_lo_lo_hi_lo,io_confOut_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_lo_hi_lo_lo = {confReg_295,confReg_294,confReg_293,confReg_292,confReg_291,confReg_290,
    confReg_289,confReg_288}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_lo_lo_hi_lo = {confReg_303,confReg_302,confReg_301,confReg_300,confReg_299,confReg_298,
    confReg_297,confReg_296,io_confOut_hi_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_lo_hi_hi_lo = {confReg_311,confReg_310,confReg_309,confReg_308,confReg_307,confReg_306,
    confReg_305,confReg_304}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_lo_lo_hi = {confReg_319,confReg_318,confReg_317,confReg_316,confReg_315,confReg_314,
    confReg_313,confReg_312,io_confOut_hi_lo_lo_hi_hi_lo,io_confOut_hi_lo_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_hi_lo_lo_lo = {confReg_327,confReg_326,confReg_325,confReg_324,confReg_323,confReg_322,
    confReg_321,confReg_320}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_lo_hi_lo_lo = {confReg_335,confReg_334,confReg_333,confReg_332,confReg_331,confReg_330,
    confReg_329,confReg_328,io_confOut_hi_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_hi_lo_hi_lo = {confReg_343,confReg_342,confReg_341,confReg_340,confReg_339,confReg_338,
    confReg_337,confReg_336}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_lo_hi_lo = {confReg_351,confReg_350,confReg_349,confReg_348,confReg_347,confReg_346,
    confReg_345,confReg_344,io_confOut_hi_lo_hi_lo_hi_lo,io_confOut_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_hi_hi_lo_lo = {confReg_359,confReg_358,confReg_357,confReg_356,confReg_355,confReg_354,
    confReg_353,confReg_352}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_lo_hi_hi_lo = {confReg_367,confReg_366,confReg_365,confReg_364,confReg_363,confReg_362,
    confReg_361,confReg_360,io_confOut_hi_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_hi_hi_hi_lo = {confReg_375,confReg_374,confReg_373,confReg_372,confReg_371,confReg_370,
    confReg_369,confReg_368}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_lo_hi_hi = {confReg_383,confReg_382,confReg_381,confReg_380,confReg_379,confReg_378,
    confReg_377,confReg_376,io_confOut_hi_lo_hi_hi_hi_lo,io_confOut_hi_lo_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_lo_lo_lo_lo = {confReg_391,confReg_390,confReg_389,confReg_388,confReg_387,confReg_386,
    confReg_385,confReg_384}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_hi_lo_lo_lo = {confReg_399,confReg_398,confReg_397,confReg_396,confReg_395,confReg_394,
    confReg_393,confReg_392,io_confOut_hi_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_lo_lo_hi_lo = {confReg_407,confReg_406,confReg_405,confReg_404,confReg_403,confReg_402,
    confReg_401,confReg_400}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_hi_lo_lo = {confReg_415,confReg_414,confReg_413,confReg_412,confReg_411,confReg_410,
    confReg_409,confReg_408,io_confOut_hi_hi_lo_lo_hi_lo,io_confOut_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_lo_hi_lo_lo = {confReg_423,confReg_422,confReg_421,confReg_420,confReg_419,confReg_418,
    confReg_417,confReg_416}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_hi_lo_hi_lo = {confReg_431,confReg_430,confReg_429,confReg_428,confReg_427,confReg_426,
    confReg_425,confReg_424,io_confOut_hi_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_lo_hi_hi_lo = {confReg_439,confReg_438,confReg_437,confReg_436,confReg_435,confReg_434,
    confReg_433,confReg_432}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_hi_lo_hi = {confReg_447,confReg_446,confReg_445,confReg_444,confReg_443,confReg_442,
    confReg_441,confReg_440,io_confOut_hi_hi_lo_hi_hi_lo,io_confOut_hi_hi_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_hi_lo_lo_lo = {confReg_455,confReg_454,confReg_453,confReg_452,confReg_451,confReg_450,
    confReg_449,confReg_448}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_hi_hi_lo_lo = {confReg_463,confReg_462,confReg_461,confReg_460,confReg_459,confReg_458,
    confReg_457,confReg_456,io_confOut_hi_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_hi_lo_hi_lo = {confReg_471,confReg_470,confReg_469,confReg_468,confReg_467,confReg_466,
    confReg_465,confReg_464}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_hi_hi_lo = {confReg_479,confReg_478,confReg_477,confReg_476,confReg_475,confReg_474,
    confReg_473,confReg_472,io_confOut_hi_hi_hi_lo_hi_lo,io_confOut_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_hi_hi_lo_lo = {confReg_487,confReg_486,confReg_485,confReg_484,confReg_483,confReg_482,
    confReg_481,confReg_480}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_hi_hi_hi_lo = {confReg_495,confReg_494,confReg_493,confReg_492,confReg_491,confReg_490,
    confReg_489,confReg_488,io_confOut_hi_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_hi_hi_hi_lo = {confReg_503,confReg_502,confReg_501,confReg_500,confReg_499,confReg_498,
    confReg_497,confReg_496}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_hi_hi_hi = {confReg_511,confReg_510,confReg_509,confReg_508,confReg_507,confReg_506,
    confReg_505,confReg_504,io_confOut_hi_hi_hi_hi_hi_lo,io_confOut_hi_hi_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [255:0] io_confOut_hi = {io_confOut_hi_hi_hi_hi,io_confOut_hi_hi_hi_lo,io_confOut_hi_hi_lo_hi,
    io_confOut_hi_hi_lo_lo,io_confOut_hi_lo_hi_hi,io_confOut_hi_lo_hi_lo,io_confOut_hi_lo_lo_hi,io_confOut_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  assign ioBundle_confOut = {io_confOut_hi,io_confOut_lo}; // @[ScanConf.scala 48:25]
  assign ioBundle_scan_out = {io_scan_out_hi,io_scan_out_lo}; // @[ScanConf.scala 46:47]
  always @(posedge clock) begin
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_0 <= confReg_8; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_1 <= confReg_9; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_2 <= confReg_10; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_3 <= confReg_11; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_4 <= confReg_12; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_5 <= confReg_13; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_6 <= confReg_14; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_7 <= confReg_15; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_8 <= confReg_16; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_9 <= confReg_17; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_10 <= confReg_18; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_11 <= confReg_19; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_12 <= confReg_20; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_13 <= confReg_21; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_14 <= confReg_22; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_15 <= confReg_23; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_16 <= confReg_24; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_17 <= confReg_25; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_18 <= confReg_26; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_19 <= confReg_27; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_20 <= confReg_28; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_21 <= confReg_29; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_22 <= confReg_30; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_23 <= confReg_31; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_24 <= confReg_32; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_25 <= confReg_33; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_26 <= confReg_34; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_27 <= confReg_35; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_28 <= confReg_36; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_29 <= confReg_37; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_30 <= confReg_38; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_31 <= confReg_39; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_32 <= confReg_40; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_33 <= confReg_41; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_34 <= confReg_42; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_35 <= confReg_43; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_36 <= confReg_44; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_37 <= confReg_45; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_38 <= confReg_46; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_39 <= confReg_47; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_40 <= confReg_48; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_41 <= confReg_49; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_42 <= confReg_50; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_43 <= confReg_51; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_44 <= confReg_52; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_45 <= confReg_53; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_46 <= confReg_54; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_47 <= confReg_55; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_48 <= confReg_56; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_49 <= confReg_57; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_50 <= confReg_58; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_51 <= confReg_59; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_52 <= confReg_60; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_53 <= confReg_61; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_54 <= confReg_62; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_55 <= confReg_63; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_56 <= confReg_64; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_57 <= confReg_65; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_58 <= confReg_66; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_59 <= confReg_67; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_60 <= confReg_68; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_61 <= confReg_69; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_62 <= confReg_70; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_63 <= confReg_71; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_64 <= confReg_72; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_65 <= confReg_73; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_66 <= confReg_74; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_67 <= confReg_75; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_68 <= confReg_76; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_69 <= confReg_77; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_70 <= confReg_78; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_71 <= confReg_79; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_72 <= confReg_80; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_73 <= confReg_81; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_74 <= confReg_82; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_75 <= confReg_83; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_76 <= confReg_84; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_77 <= confReg_85; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_78 <= confReg_86; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_79 <= confReg_87; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_80 <= confReg_88; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_81 <= confReg_89; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_82 <= confReg_90; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_83 <= confReg_91; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_84 <= confReg_92; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_85 <= confReg_93; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_86 <= confReg_94; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_87 <= confReg_95; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_88 <= confReg_96; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_89 <= confReg_97; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_90 <= confReg_98; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_91 <= confReg_99; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_92 <= confReg_100; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_93 <= confReg_101; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_94 <= confReg_102; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_95 <= confReg_103; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_96 <= confReg_104; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_97 <= confReg_105; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_98 <= confReg_106; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_99 <= confReg_107; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_100 <= confReg_108; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_101 <= confReg_109; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_102 <= confReg_110; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_103 <= confReg_111; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_104 <= confReg_112; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_105 <= confReg_113; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_106 <= confReg_114; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_107 <= confReg_115; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_108 <= confReg_116; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_109 <= confReg_117; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_110 <= confReg_118; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_111 <= confReg_119; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_112 <= confReg_120; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_113 <= confReg_121; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_114 <= confReg_122; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_115 <= confReg_123; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_116 <= confReg_124; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_117 <= confReg_125; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_118 <= confReg_126; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_119 <= confReg_127; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_120 <= confReg_128; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_121 <= confReg_129; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_122 <= confReg_130; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_123 <= confReg_131; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_124 <= confReg_132; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_125 <= confReg_133; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_126 <= confReg_134; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_127 <= confReg_135; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_128 <= confReg_136; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_129 <= confReg_137; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_130 <= confReg_138; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_131 <= confReg_139; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_132 <= confReg_140; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_133 <= confReg_141; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_134 <= confReg_142; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_135 <= confReg_143; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_136 <= confReg_144; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_137 <= confReg_145; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_138 <= confReg_146; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_139 <= confReg_147; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_140 <= confReg_148; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_141 <= confReg_149; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_142 <= confReg_150; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_143 <= confReg_151; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_144 <= confReg_152; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_145 <= confReg_153; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_146 <= confReg_154; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_147 <= confReg_155; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_148 <= confReg_156; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_149 <= confReg_157; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_150 <= confReg_158; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_151 <= confReg_159; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_152 <= confReg_160; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_153 <= confReg_161; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_154 <= confReg_162; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_155 <= confReg_163; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_156 <= confReg_164; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_157 <= confReg_165; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_158 <= confReg_166; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_159 <= confReg_167; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_160 <= confReg_168; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_161 <= confReg_169; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_162 <= confReg_170; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_163 <= confReg_171; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_164 <= confReg_172; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_165 <= confReg_173; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_166 <= confReg_174; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_167 <= confReg_175; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_168 <= confReg_176; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_169 <= confReg_177; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_170 <= confReg_178; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_171 <= confReg_179; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_172 <= confReg_180; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_173 <= confReg_181; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_174 <= confReg_182; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_175 <= confReg_183; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_176 <= confReg_184; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_177 <= confReg_185; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_178 <= confReg_186; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_179 <= confReg_187; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_180 <= confReg_188; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_181 <= confReg_189; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_182 <= confReg_190; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_183 <= confReg_191; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_184 <= confReg_192; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_185 <= confReg_193; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_186 <= confReg_194; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_187 <= confReg_195; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_188 <= confReg_196; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_189 <= confReg_197; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_190 <= confReg_198; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_191 <= confReg_199; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_192 <= confReg_200; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_193 <= confReg_201; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_194 <= confReg_202; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_195 <= confReg_203; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_196 <= confReg_204; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_197 <= confReg_205; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_198 <= confReg_206; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_199 <= confReg_207; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_200 <= confReg_208; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_201 <= confReg_209; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_202 <= confReg_210; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_203 <= confReg_211; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_204 <= confReg_212; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_205 <= confReg_213; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_206 <= confReg_214; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_207 <= confReg_215; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_208 <= confReg_216; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_209 <= confReg_217; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_210 <= confReg_218; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_211 <= confReg_219; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_212 <= confReg_220; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_213 <= confReg_221; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_214 <= confReg_222; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_215 <= confReg_223; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_216 <= confReg_224; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_217 <= confReg_225; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_218 <= confReg_226; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_219 <= confReg_227; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_220 <= confReg_228; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_221 <= confReg_229; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_222 <= confReg_230; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_223 <= confReg_231; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_224 <= confReg_232; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_225 <= confReg_233; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_226 <= confReg_234; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_227 <= confReg_235; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_228 <= confReg_236; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_229 <= confReg_237; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_230 <= confReg_238; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_231 <= confReg_239; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_232 <= confReg_240; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_233 <= confReg_241; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_234 <= confReg_242; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_235 <= confReg_243; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_236 <= confReg_244; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_237 <= confReg_245; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_238 <= confReg_246; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_239 <= confReg_247; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_240 <= confReg_248; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_241 <= confReg_249; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_242 <= confReg_250; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_243 <= confReg_251; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_244 <= confReg_252; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_245 <= confReg_253; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_246 <= confReg_254; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_247 <= confReg_255; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_248 <= confReg_256; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_249 <= confReg_257; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_250 <= confReg_258; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_251 <= confReg_259; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_252 <= confReg_260; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_253 <= confReg_261; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_254 <= confReg_262; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_255 <= confReg_263; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_256 <= confReg_264; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_257 <= confReg_265; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_258 <= confReg_266; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_259 <= confReg_267; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_260 <= confReg_268; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_261 <= confReg_269; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_262 <= confReg_270; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_263 <= confReg_271; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_264 <= confReg_272; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_265 <= confReg_273; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_266 <= confReg_274; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_267 <= confReg_275; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_268 <= confReg_276; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_269 <= confReg_277; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_270 <= confReg_278; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_271 <= confReg_279; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_272 <= confReg_280; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_273 <= confReg_281; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_274 <= confReg_282; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_275 <= confReg_283; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_276 <= confReg_284; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_277 <= confReg_285; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_278 <= confReg_286; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_279 <= confReg_287; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_280 <= confReg_288; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_281 <= confReg_289; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_282 <= confReg_290; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_283 <= confReg_291; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_284 <= confReg_292; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_285 <= confReg_293; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_286 <= confReg_294; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_287 <= confReg_295; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_288 <= confReg_296; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_289 <= confReg_297; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_290 <= confReg_298; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_291 <= confReg_299; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_292 <= confReg_300; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_293 <= confReg_301; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_294 <= confReg_302; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_295 <= confReg_303; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_296 <= confReg_304; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_297 <= confReg_305; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_298 <= confReg_306; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_299 <= confReg_307; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_300 <= confReg_308; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_301 <= confReg_309; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_302 <= confReg_310; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_303 <= confReg_311; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_304 <= confReg_312; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_305 <= confReg_313; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_306 <= confReg_314; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_307 <= confReg_315; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_308 <= confReg_316; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_309 <= confReg_317; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_310 <= confReg_318; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_311 <= confReg_319; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_312 <= confReg_320; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_313 <= confReg_321; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_314 <= confReg_322; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_315 <= confReg_323; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_316 <= confReg_324; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_317 <= confReg_325; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_318 <= confReg_326; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_319 <= confReg_327; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_320 <= confReg_328; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_321 <= confReg_329; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_322 <= confReg_330; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_323 <= confReg_331; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_324 <= confReg_332; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_325 <= confReg_333; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_326 <= confReg_334; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_327 <= confReg_335; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_328 <= confReg_336; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_329 <= confReg_337; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_330 <= confReg_338; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_331 <= confReg_339; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_332 <= confReg_340; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_333 <= confReg_341; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_334 <= confReg_342; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_335 <= confReg_343; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_336 <= confReg_344; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_337 <= confReg_345; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_338 <= confReg_346; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_339 <= confReg_347; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_340 <= confReg_348; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_341 <= confReg_349; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_342 <= confReg_350; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_343 <= confReg_351; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_344 <= confReg_352; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_345 <= confReg_353; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_346 <= confReg_354; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_347 <= confReg_355; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_348 <= confReg_356; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_349 <= confReg_357; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_350 <= confReg_358; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_351 <= confReg_359; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_352 <= confReg_360; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_353 <= confReg_361; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_354 <= confReg_362; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_355 <= confReg_363; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_356 <= confReg_364; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_357 <= confReg_365; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_358 <= confReg_366; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_359 <= confReg_367; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_360 <= confReg_368; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_361 <= confReg_369; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_362 <= confReg_370; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_363 <= confReg_371; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_364 <= confReg_372; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_365 <= confReg_373; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_366 <= confReg_374; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_367 <= confReg_375; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_368 <= confReg_376; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_369 <= confReg_377; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_370 <= confReg_378; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_371 <= confReg_379; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_372 <= confReg_380; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_373 <= confReg_381; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_374 <= confReg_382; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_375 <= confReg_383; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_376 <= confReg_384; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_377 <= confReg_385; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_378 <= confReg_386; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_379 <= confReg_387; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_380 <= confReg_388; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_381 <= confReg_389; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_382 <= confReg_390; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_383 <= confReg_391; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_384 <= confReg_392; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_385 <= confReg_393; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_386 <= confReg_394; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_387 <= confReg_395; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_388 <= confReg_396; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_389 <= confReg_397; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_390 <= confReg_398; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_391 <= confReg_399; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_392 <= confReg_400; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_393 <= confReg_401; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_394 <= confReg_402; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_395 <= confReg_403; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_396 <= confReg_404; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_397 <= confReg_405; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_398 <= confReg_406; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_399 <= confReg_407; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_400 <= confReg_408; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_401 <= confReg_409; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_402 <= confReg_410; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_403 <= confReg_411; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_404 <= confReg_412; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_405 <= confReg_413; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_406 <= confReg_414; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_407 <= confReg_415; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_408 <= confReg_416; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_409 <= confReg_417; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_410 <= confReg_418; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_411 <= confReg_419; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_412 <= confReg_420; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_413 <= confReg_421; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_414 <= confReg_422; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_415 <= confReg_423; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_416 <= confReg_424; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_417 <= confReg_425; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_418 <= confReg_426; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_419 <= confReg_427; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_420 <= confReg_428; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_421 <= confReg_429; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_422 <= confReg_430; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_423 <= confReg_431; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_424 <= confReg_432; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_425 <= confReg_433; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_426 <= confReg_434; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_427 <= confReg_435; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_428 <= confReg_436; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_429 <= confReg_437; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_430 <= confReg_438; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_431 <= confReg_439; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_432 <= confReg_440; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_433 <= confReg_441; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_434 <= confReg_442; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_435 <= confReg_443; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_436 <= confReg_444; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_437 <= confReg_445; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_438 <= confReg_446; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_439 <= confReg_447; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_440 <= confReg_448; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_441 <= confReg_449; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_442 <= confReg_450; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_443 <= confReg_451; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_444 <= confReg_452; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_445 <= confReg_453; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_446 <= confReg_454; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_447 <= confReg_455; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_448 <= confReg_456; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_449 <= confReg_457; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_450 <= confReg_458; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_451 <= confReg_459; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_452 <= confReg_460; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_453 <= confReg_461; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_454 <= confReg_462; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_455 <= confReg_463; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_456 <= confReg_464; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_457 <= confReg_465; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_458 <= confReg_466; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_459 <= confReg_467; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_460 <= confReg_468; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_461 <= confReg_469; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_462 <= confReg_470; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_463 <= confReg_471; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_464 <= confReg_472; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_465 <= confReg_473; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_466 <= confReg_474; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_467 <= confReg_475; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_468 <= confReg_476; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_469 <= confReg_477; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_470 <= confReg_478; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_471 <= confReg_479; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_472 <= confReg_480; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_473 <= confReg_481; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_474 <= confReg_482; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_475 <= confReg_483; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_476 <= confReg_484; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_477 <= confReg_485; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_478 <= confReg_486; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_479 <= confReg_487; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_480 <= confReg_488; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_481 <= confReg_489; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_482 <= confReg_490; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_483 <= confReg_491; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_484 <= confReg_492; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_485 <= confReg_493; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_486 <= confReg_494; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_487 <= confReg_495; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_488 <= confReg_496; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_489 <= confReg_497; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_490 <= confReg_498; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_491 <= confReg_499; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_492 <= confReg_500; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_493 <= confReg_501; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_494 <= confReg_502; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_495 <= confReg_503; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_496 <= confReg_504; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_497 <= confReg_505; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_498 <= confReg_506; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_499 <= confReg_507; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_500 <= confReg_508; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_501 <= confReg_509; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_502 <= confReg_510; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_503 <= confReg_511; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_504 <= ioBundle_scan_in[0]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_505 <= ioBundle_scan_in[1]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_506 <= ioBundle_scan_in[2]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_507 <= ioBundle_scan_in[3]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_508 <= ioBundle_scan_in[4]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_509 <= ioBundle_scan_in[5]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_510 <= ioBundle_scan_in[6]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_511 <= ioBundle_scan_in[7]; // @[ScanConf.scala 38:72]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  confReg_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  confReg_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  confReg_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  confReg_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  confReg_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  confReg_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  confReg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  confReg_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  confReg_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  confReg_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  confReg_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  confReg_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  confReg_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  confReg_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  confReg_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  confReg_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  confReg_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  confReg_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  confReg_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  confReg_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  confReg_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  confReg_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  confReg_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  confReg_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  confReg_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  confReg_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  confReg_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  confReg_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  confReg_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  confReg_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  confReg_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  confReg_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  confReg_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  confReg_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  confReg_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  confReg_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  confReg_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  confReg_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  confReg_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  confReg_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  confReg_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  confReg_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  confReg_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  confReg_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  confReg_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  confReg_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  confReg_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  confReg_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  confReg_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  confReg_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  confReg_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  confReg_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  confReg_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  confReg_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  confReg_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  confReg_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  confReg_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  confReg_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  confReg_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  confReg_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  confReg_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  confReg_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  confReg_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  confReg_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  confReg_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  confReg_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  confReg_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  confReg_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  confReg_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  confReg_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  confReg_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  confReg_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  confReg_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  confReg_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  confReg_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  confReg_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  confReg_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  confReg_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  confReg_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  confReg_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  confReg_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  confReg_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  confReg_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  confReg_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  confReg_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  confReg_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  confReg_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  confReg_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  confReg_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  confReg_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  confReg_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  confReg_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  confReg_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  confReg_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  confReg_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  confReg_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  confReg_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  confReg_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  confReg_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  confReg_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  confReg_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  confReg_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  confReg_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  confReg_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  confReg_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  confReg_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  confReg_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  confReg_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  confReg_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  confReg_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  confReg_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  confReg_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  confReg_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  confReg_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  confReg_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  confReg_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  confReg_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  confReg_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  confReg_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  confReg_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  confReg_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  confReg_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  confReg_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  confReg_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  confReg_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  confReg_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  confReg_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  confReg_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  confReg_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  confReg_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  confReg_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  confReg_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  confReg_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  confReg_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  confReg_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  confReg_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  confReg_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  confReg_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  confReg_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  confReg_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  confReg_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  confReg_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  confReg_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  confReg_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  confReg_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  confReg_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  confReg_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  confReg_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  confReg_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  confReg_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  confReg_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  confReg_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  confReg_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  confReg_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  confReg_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  confReg_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  confReg_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  confReg_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  confReg_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  confReg_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  confReg_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  confReg_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  confReg_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  confReg_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  confReg_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  confReg_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  confReg_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  confReg_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  confReg_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  confReg_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  confReg_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  confReg_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  confReg_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  confReg_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  confReg_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  confReg_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  confReg_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  confReg_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  confReg_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  confReg_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  confReg_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  confReg_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  confReg_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  confReg_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  confReg_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  confReg_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  confReg_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  confReg_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  confReg_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  confReg_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  confReg_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  confReg_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  confReg_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  confReg_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  confReg_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  confReg_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  confReg_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  confReg_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  confReg_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  confReg_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  confReg_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  confReg_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  confReg_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  confReg_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  confReg_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  confReg_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  confReg_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  confReg_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  confReg_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  confReg_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  confReg_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  confReg_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  confReg_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  confReg_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  confReg_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  confReg_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  confReg_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  confReg_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  confReg_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  confReg_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  confReg_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  confReg_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  confReg_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  confReg_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  confReg_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  confReg_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  confReg_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  confReg_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  confReg_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  confReg_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  confReg_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  confReg_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  confReg_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  confReg_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  confReg_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  confReg_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  confReg_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  confReg_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  confReg_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  confReg_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  confReg_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  confReg_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  confReg_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  confReg_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  confReg_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  confReg_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  confReg_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  confReg_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  confReg_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  confReg_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  confReg_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  confReg_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  confReg_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  confReg_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  confReg_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  confReg_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  confReg_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  confReg_257 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  confReg_258 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  confReg_259 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  confReg_260 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  confReg_261 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  confReg_262 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  confReg_263 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  confReg_264 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  confReg_265 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  confReg_266 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  confReg_267 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  confReg_268 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  confReg_269 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  confReg_270 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  confReg_271 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  confReg_272 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  confReg_273 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  confReg_274 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  confReg_275 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  confReg_276 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  confReg_277 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  confReg_278 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  confReg_279 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  confReg_280 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  confReg_281 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  confReg_282 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  confReg_283 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  confReg_284 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  confReg_285 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  confReg_286 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  confReg_287 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  confReg_288 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  confReg_289 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  confReg_290 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  confReg_291 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  confReg_292 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  confReg_293 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  confReg_294 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  confReg_295 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  confReg_296 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  confReg_297 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  confReg_298 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  confReg_299 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  confReg_300 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  confReg_301 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  confReg_302 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  confReg_303 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  confReg_304 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  confReg_305 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  confReg_306 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  confReg_307 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  confReg_308 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  confReg_309 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  confReg_310 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  confReg_311 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  confReg_312 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  confReg_313 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  confReg_314 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  confReg_315 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  confReg_316 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  confReg_317 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  confReg_318 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  confReg_319 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  confReg_320 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  confReg_321 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  confReg_322 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  confReg_323 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  confReg_324 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  confReg_325 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  confReg_326 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  confReg_327 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  confReg_328 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  confReg_329 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  confReg_330 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  confReg_331 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  confReg_332 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  confReg_333 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  confReg_334 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  confReg_335 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  confReg_336 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  confReg_337 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  confReg_338 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  confReg_339 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  confReg_340 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  confReg_341 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  confReg_342 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  confReg_343 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  confReg_344 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  confReg_345 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  confReg_346 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  confReg_347 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  confReg_348 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  confReg_349 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  confReg_350 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  confReg_351 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  confReg_352 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  confReg_353 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  confReg_354 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  confReg_355 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  confReg_356 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  confReg_357 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  confReg_358 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  confReg_359 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  confReg_360 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  confReg_361 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  confReg_362 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  confReg_363 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  confReg_364 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  confReg_365 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  confReg_366 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  confReg_367 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  confReg_368 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  confReg_369 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  confReg_370 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  confReg_371 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  confReg_372 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  confReg_373 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  confReg_374 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  confReg_375 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  confReg_376 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  confReg_377 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  confReg_378 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  confReg_379 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  confReg_380 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  confReg_381 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  confReg_382 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  confReg_383 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  confReg_384 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  confReg_385 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  confReg_386 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  confReg_387 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  confReg_388 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  confReg_389 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  confReg_390 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  confReg_391 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  confReg_392 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  confReg_393 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  confReg_394 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  confReg_395 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  confReg_396 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  confReg_397 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  confReg_398 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  confReg_399 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  confReg_400 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  confReg_401 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  confReg_402 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  confReg_403 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  confReg_404 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  confReg_405 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  confReg_406 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  confReg_407 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  confReg_408 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  confReg_409 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  confReg_410 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  confReg_411 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  confReg_412 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  confReg_413 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  confReg_414 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  confReg_415 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  confReg_416 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  confReg_417 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  confReg_418 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  confReg_419 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  confReg_420 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  confReg_421 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  confReg_422 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  confReg_423 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  confReg_424 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  confReg_425 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  confReg_426 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  confReg_427 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  confReg_428 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  confReg_429 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  confReg_430 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  confReg_431 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  confReg_432 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  confReg_433 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  confReg_434 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  confReg_435 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  confReg_436 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  confReg_437 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  confReg_438 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  confReg_439 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  confReg_440 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  confReg_441 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  confReg_442 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  confReg_443 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  confReg_444 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  confReg_445 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  confReg_446 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  confReg_447 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  confReg_448 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  confReg_449 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  confReg_450 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  confReg_451 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  confReg_452 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  confReg_453 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  confReg_454 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  confReg_455 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  confReg_456 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  confReg_457 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  confReg_458 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  confReg_459 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  confReg_460 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  confReg_461 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  confReg_462 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  confReg_463 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  confReg_464 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  confReg_465 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  confReg_466 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  confReg_467 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  confReg_468 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  confReg_469 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  confReg_470 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  confReg_471 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  confReg_472 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  confReg_473 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  confReg_474 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  confReg_475 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  confReg_476 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  confReg_477 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  confReg_478 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  confReg_479 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  confReg_480 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  confReg_481 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  confReg_482 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  confReg_483 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  confReg_484 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  confReg_485 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  confReg_486 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  confReg_487 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  confReg_488 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  confReg_489 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  confReg_490 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  confReg_491 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  confReg_492 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  confReg_493 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  confReg_494 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  confReg_495 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  confReg_496 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  confReg_497 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  confReg_498 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  confReg_499 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  confReg_500 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  confReg_501 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  confReg_502 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  confReg_503 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  confReg_504 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  confReg_505 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  confReg_506 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  confReg_507 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  confReg_508 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  confReg_509 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  confReg_510 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  confReg_511 = _RAND_511[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MuxNInput_10_SCAOptCB(
  input  [9:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_cnstClk,
  input        io_arst
);
  wire [15:0] OPinMux_in; // @[MuxListTest.scala 43:28]
  wire [3:0] OPinMux_sel; // @[MuxListTest.scala 43:28]
  wire  OPinMux_o; // @[MuxListTest.scala 43:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux16C OPinMux ( // @[MuxListTest.scala 43:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{6'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_12_SCAOptCB(
  input  [11:0] io_in,
  input  [3:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [15:0] OPinMux_in; // @[MuxListTest.scala 43:28]
  wire [3:0] OPinMux_sel; // @[MuxListTest.scala 43:28]
  wire  OPinMux_o; // @[MuxListTest.scala 43:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux16C OPinMux ( // @[MuxListTest.scala 43:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{4'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_16_SCAOptCB(
  input  [15:0] io_in,
  input  [4:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [31:0] OPinMux_in; // @[MuxListTest.scala 44:28]
  wire [4:0] OPinMux_sel; // @[MuxListTest.scala 44:28]
  wire  OPinMux_o; // @[MuxListTest.scala 44:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux32C OPinMux ( // @[MuxListTest.scala 44:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{16'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_14_SCAOptCB(
  input  [13:0] io_in,
  input  [3:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [15:0] OPinMux_in; // @[MuxListTest.scala 43:28]
  wire [3:0] OPinMux_sel; // @[MuxListTest.scala 43:28]
  wire  OPinMux_o; // @[MuxListTest.scala 43:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux16C OPinMux ( // @[MuxListTest.scala 43:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{2'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_8_SCAOptCB(
  input  [7:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_cnstClk,
  input        io_arst
);
  wire [15:0] OPinMux_in; // @[MuxListTest.scala 43:28]
  wire [3:0] OPinMux_sel; // @[MuxListTest.scala 43:28]
  wire  OPinMux_o; // @[MuxListTest.scala 43:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux16C OPinMux ( // @[MuxListTest.scala 43:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{8'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_1_SCAOptCB(
  input   io_in,
  input   io_config,
  output  io_out,
  input   io_loopBreak,
  input   io_cnstClk,
  input   io_arst
);
  wire [1:0] OPinMux_in; // @[MuxListTest.scala 40:28]
  wire  OPinMux_sel; // @[MuxListTest.scala 40:28]
  wire  OPinMux_o; // @[MuxListTest.scala 40:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux2C OPinMux ( // @[MuxListTest.scala 40:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{1'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_O3_C6_SCAOptSB(
  input  [8:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{5'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in[8:3]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O4_C5_SCAOptSB(
  input  [8:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{4'd0}, io_in[3:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in[8:4]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O4_C6_SCAOptSB(
  input  [9:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{4'd0}, io_in[3:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in[9:4]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O0_C6_SCAOptSB(
  input  [5:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = 8'h0; // @[MuxListTest.scala 125:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O3_C5_SCAOptSB(
  input  [7:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{5'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in[7:3]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O0_C4_SCAOptSB(
  input  [3:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = 4'h0; // @[MuxListTest.scala 125:22]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = io_in; // @[MuxListTest.scala 144:28]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O4_C7_SCAOptSB(
  input  [10:0] io_in,
  input  [3:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_ioGndBle,
  input         io_cnstClk,
  input         io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{4'd0}, io_in[3:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{1'd0}, io_in[10:4]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O3_C7_SCAOptSB(
  input  [9:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{5'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{1'd0}, io_in[9:3]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module Tile_3_3_clbalutile(
  input          clock,
  input          reset,
  input          IN_OPIN_N5807_73,
  input          IN_OPIN_N5808_74,
  input          IN_OPIN_N5809_75,
  input          IN_OPIN_N5810_76,
  input          IN_OPIN_N5811_77,
  input          IN_OPIN_N5812_78,
  input          IN_OPIN_N5813_79,
  input          IN_OPIN_N5814_80,
  input          IN_OPIN_N5823_89,
  input          IN_OPIN_N5824_90,
  input          IN_OPIN_N5825_91,
  input          IN_OPIN_N5826_92,
  input          IN_OPIN_N5827_93,
  input          IN_OPIN_N5828_94,
  input          IN_OPIN_N5829_95,
  input          IN_OPIN_N5830_96,
  input          IN_OPIN_N5831_97,
  input          IN_OPIN_N5832_98,
  input          IN_OPIN_N5833_99,
  input          IN_OPIN_N5834_100,
  input          IN_OPIN_N5835_101,
  input          IN_OPIN_N5836_102,
  input          IN_OPIN_N5837_103,
  input          IN_OPIN_N5838_104,
  input          IN_OPIN_N5839_105,
  input          IN_OPIN_N5840_106,
  input          IN_OPIN_N5841_107,
  input          IN_OPIN_N5842_108,
  input          IN_OPIN_N5843_109,
  input          IN_OPIN_N5844_110,
  input          IN_OPIN_N5845_111,
  input          IN_OPIN_N5846_112,
  input          IN_OPIN_N5847_113,
  input          IN_OPIN_N5848_114,
  input          IN_OPIN_N5849_115,
  input          IN_OPIN_N5850_116,
  input          IN_OPIN_N5851_117,
  input          IN_OPIN_N5852_118,
  input          IN_OPIN_N5853_119,
  input          IN_OPIN_N5854_120,
  input          IN_OPIN_N8011_81,
  input          IN_OPIN_N8012_82,
  input          IN_OPIN_N8013_83,
  input          IN_OPIN_N8014_84,
  input          IN_OPIN_N8015_85,
  input          IN_OPIN_N8016_86,
  input          IN_OPIN_N8017_87,
  input          IN_OPIN_N8018_88,
  input          IN_CHANX_N23992_4,
  input          IN_CHANX_N23994_6,
  input          IN_CHANX_N23995_7,
  input          IN_CHANX_N24000_12,
  input          IN_CHANX_N24002_14,
  input          IN_CHANX_N24003_15,
  input          IN_CHANX_N24008_20,
  input          IN_CHANX_N24010_22,
  input          IN_CHANX_N24011_23,
  input          IN_CHANX_N24016_28,
  input          IN_CHANX_N24018_30,
  input          IN_CHANX_N24019_31,
  input          IN_CHANX_N24024_36,
  input          IN_CHANX_N24032_44,
  input          IN_CHANX_N24040_52,
  input          IN_CHANX_N24048_60,
  input          IN_CHANX_N24056_68,
  input          IN_CHANX_N24068_0,
  input          IN_CHANX_N24069_1,
  input          IN_CHANX_N24070_8,
  input          IN_CHANX_N24071_9,
  input          IN_CHANX_N24072_16,
  input          IN_CHANX_N24073_17,
  input          IN_CHANX_N24074_24,
  input          IN_CHANX_N24075_25,
  input          IN_CHANX_N24076_32,
  input          IN_CHANX_N24077_33,
  input          IN_CHANX_N24088_76,
  input          IN_CHANX_N24090_2,
  input          IN_CHANX_N24091_3,
  input          IN_CHANX_N24092_10,
  input          IN_CHANX_N24093_11,
  input          IN_CHANX_N24094_18,
  input          IN_CHANX_N24095_19,
  input          IN_CHANX_N24096_26,
  input          IN_CHANX_N24097_27,
  input          IN_CHANX_N24098_34,
  input          IN_CHANX_N24099_35,
  input          IN_CHANX_N24100_42,
  input          IN_CHANX_N24101_43,
  input          IN_CHANX_N24102_50,
  input          IN_CHANX_N24103_51,
  input          IN_CHANX_N24104_58,
  input          IN_CHANX_N24105_59,
  input          IN_CHANX_N24106_66,
  input          IN_CHANX_N24107_67,
  input          IN_CHANX_N24108_74,
  input          IN_CHANX_N24109_75,
  input          IN_CHANX_N24113_5,
  input          IN_CHANX_N24115_13,
  input          IN_CHANX_N24117_21,
  input          IN_CHANX_N24119_29,
  input          IN_CHANX_N24121_37,
  input          IN_CHANX_N24123_45,
  input          IN_CHANX_N24125_53,
  input          IN_CHANX_N24127_61,
  input          IN_CHANX_N24129_69,
  input          IN_CHANX_N24131_77,
  input          IN_CHANY_N27118_4,
  input          IN_CHANY_N27120_6,
  input          IN_CHANY_N27121_7,
  input          IN_CHANY_N27126_12,
  input          IN_CHANY_N27128_14,
  input          IN_CHANY_N27129_15,
  input          IN_CHANY_N27134_20,
  input          IN_CHANY_N27136_22,
  input          IN_CHANY_N27137_23,
  input          IN_CHANY_N27142_28,
  input          IN_CHANY_N27144_30,
  input          IN_CHANY_N27145_31,
  input          IN_CHANY_N27150_36,
  input          IN_CHANY_N27158_44,
  input          IN_CHANY_N27166_52,
  input          IN_CHANY_N27174_60,
  input          IN_CHANY_N27182_68,
  input          IN_CHANY_N27194_0,
  input          IN_CHANY_N27195_1,
  input          IN_CHANY_N27196_8,
  input          IN_CHANY_N27197_9,
  input          IN_CHANY_N27198_16,
  input          IN_CHANY_N27199_17,
  input          IN_CHANY_N27200_24,
  input          IN_CHANY_N27201_25,
  input          IN_CHANY_N27202_32,
  input          IN_CHANY_N27203_33,
  input          IN_CHANY_N27214_76,
  input          IN_CHANY_N27216_2,
  input          IN_CHANY_N27217_3,
  input          IN_CHANY_N27218_10,
  input          IN_CHANY_N27219_11,
  input          IN_CHANY_N27220_18,
  input          IN_CHANY_N27221_19,
  input          IN_CHANY_N27222_26,
  input          IN_CHANY_N27223_27,
  input          IN_CHANY_N27224_34,
  input          IN_CHANY_N27225_35,
  input          IN_CHANY_N27226_42,
  input          IN_CHANY_N27227_43,
  input          IN_CHANY_N27228_50,
  input          IN_CHANY_N27229_51,
  input          IN_CHANY_N27230_58,
  input          IN_CHANY_N27231_59,
  input          IN_CHANY_N27232_66,
  input          IN_CHANY_N27233_67,
  input          IN_CHANY_N27234_74,
  input          IN_CHANY_N27235_75,
  input          IN_CHANY_N27236_78,
  input          IN_CHANY_N27237_79,
  input          IN_CHANY_N27239_5,
  input          IN_CHANY_N27241_13,
  input          IN_CHANY_N27243_21,
  input          IN_CHANY_N27245_29,
  input          IN_CHANY_N27247_37,
  input          IN_CHANY_N27249_45,
  input          IN_CHANY_N27251_53,
  input          IN_CHANY_N27253_61,
  input          IN_CHANY_N27255_69,
  input          IN_CHANY_N27257_77,
  output         OUT_OPIN_N5581_91,
  output         OUT_OPIN_N5603_113,
  output         OUT_OPIN_N5572_82,
  output         OUT_OPIN_N5610_120,
  output         OUT_CHANY_N27159_45,
  output         OUT_CHANX_N24009_21,
  output         OUT_OPIN_N5577_87,
  output         OUT_CHANY_N27240_12,
  output         OUT_CHANY_N27151_37,
  output         OUT_OPIN_N5600_110,
  output         OUT_OPIN_N5566_76,
  output         OUT_CHANY_N27254_68,
  output         OUT_CHANY_N27143_29,
  output         OUT_OPIN_N5595_105,
  output         OUT_CHANX_N24120_36,
  output         OUT_CHANY_N27244_28,
  output         OUT_OPIN_N5601_111,
  output         OUT_CHANY_N27242_20,
  output         OUT_CHANY_N27119_5,
  output         OUT_OPIN_N5609_119,
  output         OUT_OPIN_N5588_98,
  output         OUT_CHANX_N24126_60,
  output         OUT_OPIN_N5604_114,
  output         OUT_CHANX_N24033_45,
  output         OUT_CHANY_N27175_61,
  output         OUT_CHANY_N27250_52,
  output         OUT_CHANX_N24112_4,
  output         OUT_CHANX_N24057_69,
  output         OUT_CHANX_N24130_76,
  output         OUT_CHANY_N27252_60,
  output         OUT_OPIN_N5585_95,
  output         OUT_CHANY_N27246_36,
  output         OUT_OPIN_N5586_96,
  output         OUT_CHANX_N24041_53,
  output         OUT_OPIN_N5568_78,
  output         OUT_OPIN_N5592_102,
  output         OUT_OPIN_N5583_93,
  output         OUT_OPIN_N5605_115,
  output         OUT_OPIN_N5608_118,
  output         OUT_CHANX_N24118_28,
  output         OUT_OPIN_N5596_106,
  output         OUT_OPIN_N5571_81,
  output         OUT_OPIN_N5563_73,
  output         OUT_OPIN_N5576_86,
  output         OUT_OPIN_N5582_92,
  output         OUT_CHANX_N24128_68,
  output         OUT_OPIN_N5573_83,
  output         OUT_CHANX_N24017_29,
  output         OUT_OPIN_N5580_90,
  output         OUT_OPIN_N5606_116,
  output         OUT_CHANX_N24124_52,
  output         OUT_OPIN_N5598_108,
  output         OUT_CHANX_N24049_61,
  output         OUT_OPIN_N5589_99,
  output         OUT_OPIN_N5567_77,
  output         OUT_OPIN_N5591_101,
  output         OUT_OPIN_N5597_107,
  output         OUT_OPIN_N5569_79,
  output         OUT_CHANY_N27238_4,
  output         OUT_OPIN_N5570_80,
  output         OUT_CHANY_N27183_69,
  output         OUT_OPIN_N5593_103,
  output         OUT_OPIN_N5574_84,
  output         OUT_CHANX_N24114_12,
  output         OUT_OPIN_N5575_85,
  output         OUT_OPIN_N5599_109,
  output         OUT_OPIN_N5584_94,
  output         OUT_OPIN_N5578_88,
  output         OUT_OPIN_N5579_89,
  output         OUT_CHANX_N24025_37,
  output         OUT_OPIN_N5565_75,
  output         OUT_OPIN_N5564_74,
  output         OUT_OPIN_N5587_97,
  output         OUT_CHANY_N27215_77,
  output         OUT_OPIN_N5607_117,
  output         OUT_CHANY_N27256_76,
  output         OUT_CHANX_N23993_5,
  output         OUT_OPIN_N5594_104,
  output         OUT_CHANY_N27135_21,
  output         OUT_CHANY_N27167_53,
  output         OUT_CHANX_N24001_13,
  output         OUT_CHANY_N27127_13,
  output         OUT_OPIN_N5590_100,
  output         OUT_CHANX_N24116_20,
  output         OUT_CHANX_N24122_44,
  output         OUT_CHANY_N27248_44,
  output         OUT_OPIN_N5602_112,
  output         OUT_CHANX_N24089_77,
  output [511:0] ioConf_confOut,
  input  [7:0]   ioConf_scan_in,
  input          ioConf_scan_en,
  output [7:0]   ioConf_scan_out,
  input          ctrlSignals_gndBlkOuts,
  input          ctrlSignals_loopBreak,
  input          ctrlSignals_arst,
  input          ctrlSignals_tmrMode,
  input          ctrlSignals_confClock,
  input          ctrlSignals_constClock
);
  wire  logicBlock_IPIN_0; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_1; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_2; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_3; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_4; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_5; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_6; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_7; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_8; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_9; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_10; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_11; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_12; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_13; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_14; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_15; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_16; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_17; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_18; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_19; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_20; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_21; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_22; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_23; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_24; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_25; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_26; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_27; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_28; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_29; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_30; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_31; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_32; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_33; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_34; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_35; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_36; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_37; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_38; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_39; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_40; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_41; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_42; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_43; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_44; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_45; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_46; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_47; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_48; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_49; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_50; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_51; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_52; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_53; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_54; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_55; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_56; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_57; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_58; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_59; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_60; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_61; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_62; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_63; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_64; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_65; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_66; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_67; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_68; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_69; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_70; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_71; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_73; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_74; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_75; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_76; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_77; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_78; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_79; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_80; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_81; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_82; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_83; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_84; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_85; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_86; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_87; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_88; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_89; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_90; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_91; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_92; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_93; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_94; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_95; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_96; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_97; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_98; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_99; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_100; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_101; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_102; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_103; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_104; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_105; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_106; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_107; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_108; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_109; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_110; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_111; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_112; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_113; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_114; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_115; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_116; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_117; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_118; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_119; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_120; // @[TileFull.scala 47:37]
  wire  logicBlock_clock; // @[TileFull.scala 47:37]
  wire  logicBlock_reset; // @[TileFull.scala 47:37]
  wire [193:0] logicBlock_configBits; // @[TileFull.scala 47:37]
  wire  logicBlock_gndLBouts; // @[TileFull.scala 47:37]
  wire  configBlock_clock; // @[TileFull.scala 61:31]
  wire [511:0] configBlock_ioBundle_confOut; // @[TileFull.scala 61:31]
  wire [7:0] configBlock_ioBundle_scan_in; // @[TileFull.scala 61:31]
  wire  configBlock_ioBundle_scan_en; // @[TileFull.scala 61:31]
  wire [7:0] configBlock_ioBundle_scan_out; // @[TileFull.scala 61:31]
  wire [9:0] CBMux_IPIN0_N5490_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN0_N5490_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N5490_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N5490_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N5490_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N5490_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN1_N5491_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN1_N5491_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN1_N5491_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN1_N5491_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN1_N5491_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN1_N5491_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN2_N5492_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN2_N5492_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N5492_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N5492_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N5492_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N5492_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN3_N5493_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN3_N5493_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN3_N5493_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN3_N5493_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN3_N5493_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN3_N5493_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN4_N5494_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN4_N5494_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N5494_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N5494_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N5494_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N5494_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN5_N5495_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN5_N5495_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN5_N5495_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN5_N5495_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN5_N5495_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN5_N5495_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN6_N5496_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN6_N5496_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N5496_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N5496_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N5496_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N5496_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN7_N5497_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN7_N5497_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN7_N5497_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN7_N5497_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN7_N5497_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN7_N5497_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN8_N5498_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN8_N5498_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N5498_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N5498_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N5498_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N5498_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN9_N5499_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN9_N5499_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN9_N5499_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN9_N5499_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN9_N5499_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN9_N5499_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN10_N5500_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN10_N5500_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N5500_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N5500_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N5500_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N5500_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN11_N5501_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN11_N5501_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN11_N5501_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN11_N5501_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN11_N5501_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN11_N5501_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN12_N5502_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN12_N5502_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N5502_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N5502_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N5502_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N5502_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN13_N5503_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN13_N5503_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN13_N5503_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN13_N5503_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN13_N5503_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN13_N5503_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN14_N5504_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN14_N5504_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N5504_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N5504_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N5504_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N5504_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN15_N5505_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN15_N5505_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN15_N5505_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN15_N5505_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN15_N5505_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN15_N5505_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN16_N5506_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN16_N5506_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N5506_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N5506_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N5506_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N5506_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN17_N5507_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN17_N5507_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN17_N5507_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN17_N5507_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN17_N5507_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN17_N5507_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN18_N5508_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN18_N5508_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N5508_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N5508_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N5508_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N5508_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN19_N5509_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN19_N5509_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN19_N5509_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN19_N5509_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN19_N5509_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN19_N5509_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN20_N5510_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN20_N5510_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N5510_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N5510_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N5510_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N5510_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN21_N5511_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN21_N5511_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN21_N5511_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN21_N5511_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN21_N5511_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN21_N5511_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN22_N5512_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN22_N5512_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N5512_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N5512_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N5512_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N5512_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN23_N5513_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN23_N5513_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN23_N5513_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN23_N5513_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN23_N5513_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN23_N5513_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN24_N5514_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN24_N5514_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N5514_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N5514_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N5514_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N5514_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN25_N5515_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN25_N5515_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN25_N5515_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN25_N5515_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN25_N5515_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN25_N5515_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN26_N5516_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN26_N5516_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N5516_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N5516_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N5516_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N5516_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN27_N5517_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN27_N5517_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN27_N5517_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN27_N5517_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN27_N5517_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN27_N5517_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN28_N5518_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN28_N5518_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N5518_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N5518_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N5518_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N5518_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN29_N5519_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN29_N5519_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN29_N5519_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN29_N5519_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN29_N5519_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN29_N5519_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN30_N5520_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN30_N5520_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N5520_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N5520_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N5520_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N5520_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN31_N5521_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN31_N5521_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN31_N5521_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN31_N5521_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN31_N5521_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN31_N5521_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN32_N5522_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN32_N5522_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N5522_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N5522_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N5522_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N5522_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN33_N5523_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN33_N5523_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN33_N5523_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN33_N5523_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN33_N5523_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN33_N5523_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN34_N5524_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN34_N5524_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N5524_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N5524_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N5524_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N5524_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN35_N5525_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN35_N5525_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN35_N5525_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN35_N5525_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN35_N5525_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN35_N5525_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN36_N5526_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN36_N5526_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N5526_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N5526_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N5526_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N5526_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN37_N5527_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN37_N5527_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN37_N5527_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN37_N5527_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN37_N5527_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN37_N5527_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN38_N5528_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN38_N5528_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N5528_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N5528_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N5528_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N5528_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN39_N5529_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN39_N5529_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN39_N5529_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN39_N5529_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN39_N5529_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN39_N5529_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN40_N5530_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN40_N5530_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN40_N5530_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN40_N5530_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN40_N5530_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN40_N5530_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN41_N5531_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN41_N5531_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN41_N5531_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN41_N5531_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN41_N5531_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN41_N5531_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN42_N5532_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN42_N5532_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN42_N5532_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN42_N5532_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN42_N5532_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN42_N5532_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN43_N5533_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN43_N5533_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN43_N5533_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN43_N5533_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN43_N5533_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN43_N5533_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN44_N5534_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN44_N5534_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN44_N5534_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN44_N5534_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN44_N5534_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN44_N5534_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN45_N5535_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN45_N5535_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN45_N5535_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN45_N5535_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN45_N5535_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN45_N5535_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN46_N5536_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN46_N5536_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN46_N5536_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN46_N5536_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN46_N5536_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN46_N5536_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN47_N5537_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN47_N5537_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN47_N5537_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN47_N5537_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN47_N5537_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN47_N5537_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN48_N5538_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN48_N5538_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN48_N5538_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN48_N5538_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN48_N5538_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN48_N5538_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN49_N5539_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN49_N5539_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN49_N5539_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN49_N5539_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN49_N5539_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN49_N5539_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN50_N5540_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN50_N5540_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN50_N5540_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN50_N5540_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN50_N5540_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN50_N5540_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN51_N5541_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN51_N5541_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN51_N5541_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN51_N5541_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN51_N5541_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN51_N5541_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN52_N5542_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN52_N5542_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN52_N5542_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN52_N5542_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN52_N5542_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN52_N5542_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN53_N5543_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN53_N5543_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN53_N5543_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN53_N5543_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN53_N5543_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN53_N5543_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN54_N5544_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN54_N5544_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN54_N5544_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN54_N5544_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN54_N5544_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN54_N5544_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN55_N5545_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN55_N5545_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN55_N5545_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN55_N5545_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN55_N5545_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN55_N5545_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN56_N5546_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN56_N5546_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN56_N5546_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN56_N5546_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN56_N5546_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN56_N5546_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN57_N5547_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN57_N5547_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN57_N5547_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN57_N5547_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN57_N5547_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN57_N5547_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN58_N5548_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN58_N5548_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN58_N5548_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN58_N5548_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN58_N5548_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN58_N5548_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN59_N5549_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN59_N5549_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN59_N5549_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN59_N5549_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN59_N5549_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN59_N5549_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN60_N5550_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN60_N5550_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN60_N5550_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN60_N5550_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN60_N5550_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN60_N5550_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN61_N5551_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN61_N5551_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN61_N5551_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN61_N5551_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN61_N5551_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN61_N5551_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN62_N5552_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN62_N5552_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN62_N5552_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN62_N5552_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN62_N5552_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN62_N5552_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN63_N5553_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN63_N5553_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN63_N5553_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN63_N5553_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN63_N5553_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN63_N5553_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN64_N5554_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN64_N5554_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN64_N5554_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN64_N5554_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN64_N5554_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN64_N5554_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN65_N5555_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN65_N5555_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN65_N5555_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN65_N5555_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN65_N5555_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN65_N5555_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN66_N5556_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN66_N5556_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN66_N5556_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN66_N5556_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN66_N5556_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN66_N5556_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN67_N5557_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN67_N5557_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN67_N5557_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN67_N5557_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN67_N5557_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN67_N5557_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN68_N5558_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN68_N5558_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN68_N5558_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN68_N5558_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN68_N5558_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN68_N5558_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN69_N5559_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN69_N5559_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN69_N5559_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN69_N5559_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN69_N5559_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN69_N5559_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN70_N5560_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN70_N5560_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN70_N5560_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN70_N5560_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN70_N5560_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN70_N5560_io_arst; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN71_N5561_io_in; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN71_N5561_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN71_N5561_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN71_N5561_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN71_N5561_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN71_N5561_io_arst; // @[TileFull.scala 97:27]
  wire [8:0] SBMux_C5_N23993_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C5_N23993_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N23993_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N23993_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N23993_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N23993_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N23993_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C13_N24001_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C13_N24001_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N24001_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N24001_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N24001_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N24001_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N24001_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C21_N24009_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C21_N24009_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N24009_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N24009_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N24009_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N24009_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N24009_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C29_N24017_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C29_N24017_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N24017_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N24017_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N24017_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N24017_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N24017_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C37_N24025_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C37_N24025_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N24025_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N24025_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N24025_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N24025_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N24025_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C45_N24033_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C45_N24033_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N24033_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N24033_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N24033_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N24033_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N24033_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C53_N24041_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C53_N24041_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N24041_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N24041_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N24041_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N24041_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N24041_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [9:0] SBMux_C61_N24049_O_4_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C61_N24049_O_4_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N24049_O_4_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N24049_O_4_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N24049_O_4_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N24049_O_4_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N24049_O_4_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C69_N24057_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C69_N24057_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N24057_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N24057_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N24057_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N24057_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N24057_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [5:0] SBMux_C77_N24089_O_0_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C77_N24089_O_0_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24089_O_0_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24089_O_0_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24089_O_0_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24089_O_0_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24089_O_0_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C4_N24112_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C4_N24112_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N24112_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N24112_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N24112_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N24112_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N24112_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C12_N24114_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C12_N24114_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N24114_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N24114_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N24114_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N24114_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N24114_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C20_N24116_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C20_N24116_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N24116_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N24116_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N24116_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N24116_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N24116_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C28_N24118_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C28_N24118_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N24118_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N24118_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N24118_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N24118_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N24118_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C36_N24120_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C36_N24120_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N24120_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N24120_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N24120_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N24120_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N24120_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C44_N24122_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C44_N24122_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N24122_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N24122_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N24122_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N24122_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N24122_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C52_N24124_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C52_N24124_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N24124_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N24124_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N24124_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N24124_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N24124_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C60_N24126_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C60_N24126_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N24126_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N24126_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N24126_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N24126_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N24126_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C68_N24128_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C68_N24128_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N24128_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N24128_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N24128_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N24128_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N24128_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C76_N24130_O_0_C_4_io_in; // @[TileFull.scala 134:27]
  wire [2:0] SBMux_C76_N24130_O_0_C_4_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N24130_O_0_C_4_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N24130_O_0_C_4_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N24130_O_0_C_4_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N24130_O_0_C_4_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N24130_O_0_C_4_io_arst; // @[TileFull.scala 134:27]
  wire [9:0] SBMux_C5_N27119_O_4_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C5_N27119_O_4_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N27119_O_4_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N27119_O_4_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N27119_O_4_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N27119_O_4_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N27119_O_4_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C13_N27127_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C13_N27127_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N27127_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N27127_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N27127_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N27127_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N27127_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C21_N27135_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C21_N27135_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N27135_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N27135_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N27135_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N27135_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N27135_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C29_N27143_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C29_N27143_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N27143_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N27143_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N27143_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N27143_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N27143_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C37_N27151_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C37_N27151_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N27151_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N27151_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N27151_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N27151_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N27151_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C45_N27159_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C45_N27159_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N27159_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N27159_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N27159_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N27159_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N27159_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C53_N27167_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C53_N27167_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N27167_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N27167_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N27167_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N27167_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N27167_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C61_N27175_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C61_N27175_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N27175_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N27175_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N27175_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N27175_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N27175_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C69_N27183_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C69_N27183_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N27183_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N27183_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N27183_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N27183_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N27183_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C77_N27215_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C77_N27215_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N27215_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N27215_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N27215_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N27215_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N27215_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [10:0] SBMux_C4_N27238_O_4_C_7_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C4_N27238_O_4_C_7_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N27238_O_4_C_7_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N27238_O_4_C_7_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N27238_O_4_C_7_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N27238_O_4_C_7_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N27238_O_4_C_7_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C12_N27240_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C12_N27240_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N27240_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N27240_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N27240_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N27240_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N27240_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C20_N27242_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C20_N27242_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N27242_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N27242_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N27242_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N27242_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N27242_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C28_N27244_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C28_N27244_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N27244_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N27244_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N27244_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N27244_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N27244_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C36_N27246_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C36_N27246_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N27246_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N27246_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N27246_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N27246_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N27246_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C44_N27248_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C44_N27248_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N27248_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N27248_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N27248_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N27248_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N27248_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C52_N27250_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C52_N27250_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N27250_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N27250_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N27250_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N27250_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N27250_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [9:0] SBMux_C60_N27252_O_4_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C60_N27252_O_4_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N27252_O_4_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N27252_O_4_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N27252_O_4_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N27252_O_4_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N27252_O_4_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [9:0] SBMux_C68_N27254_O_4_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C68_N27254_O_4_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N27254_O_4_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N27254_O_4_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N27254_O_4_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N27254_O_4_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N27254_O_4_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [9:0] SBMux_C76_N27256_O_3_C_7_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C76_N27256_O_3_C_7_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N27256_O_3_C_7_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N27256_O_3_C_7_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N27256_O_3_C_7_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N27256_O_3_C_7_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N27256_O_3_C_7_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] CBMux_IPIN0_N5490_io_in_lo = {IN_CHANY_N27198_16,IN_CHANY_N27129_15,IN_CHANY_N27128_14,IN_CHANY_N27121_7,
    IN_CHANY_N27120_6}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN0_N5490_io_in_hi = {IN_CHANY_N27237_79,IN_CHANY_N27236_78,IN_CHANY_N27223_27,IN_CHANY_N27222_26,
    IN_CHANY_N27199_17}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN1_N5491_io_in_WIRE_1 = SBMux_C29_N27143_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [5:0] CBMux_IPIN1_N5491_io_in_lo = {IN_CHANY_N27197_9,IN_CHANY_N27196_8,IN_CHANY_N27195_1,IN_CHANY_N27194_0,
    _CBMux_IPIN1_N5491_io_in_WIRE_1,IN_CHANY_N27142_28}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN1_N5491_io_in_WIRE_7 = SBMux_C77_N27215_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [5:0] CBMux_IPIN1_N5491_io_in_hi = {IN_CHANY_N27233_67,IN_CHANY_N27232_66,IN_CHANY_N27221_19,IN_CHANY_N27220_18,
    _CBMux_IPIN1_N5491_io_in_WIRE_7,IN_CHANY_N27214_76}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN2_N5492_io_in_WIRE_1 = SBMux_C21_N27135_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire [5:0] CBMux_IPIN2_N5492_io_in_lo = {IN_CHANY_N27217_3,IN_CHANY_N27216_2,_CBMux_IPIN1_N5491_io_in_WIRE_7,
    IN_CHANY_N27214_76,_CBMux_IPIN2_N5492_io_in_WIRE_1,IN_CHANY_N27134_20}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN2_N5492_io_in_hi = {IN_CHANY_N27231_59,IN_CHANY_N27230_58,IN_CHANY_N27225_35,IN_CHANY_N27224_34,
    IN_CHANY_N27219_11,IN_CHANY_N27218_10}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN3_N5493_io_in_WIRE_1 = SBMux_C5_N27119_O_4_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN3_N5493_io_in_WIRE_3 = SBMux_C13_N27127_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN3_N5493_io_in_WIRE_7 = SBMux_C37_N27151_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [7:0] CBMux_IPIN3_N5493_io_in_lo = {_CBMux_IPIN3_N5493_io_in_WIRE_7,IN_CHANY_N27150_36,IN_CHANY_N27145_31,
    IN_CHANY_N27144_30,_CBMux_IPIN3_N5493_io_in_WIRE_3,IN_CHANY_N27126_12,_CBMux_IPIN3_N5493_io_in_WIRE_1,
    IN_CHANY_N27118_4}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN3_N5493_io_in_hi = {IN_CHANY_N27237_79,IN_CHANY_N27236_78,IN_CHANY_N27235_75,IN_CHANY_N27234_74,
    IN_CHANY_N27229_51,IN_CHANY_N27228_50,IN_CHANY_N27227_43,IN_CHANY_N27226_42}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN4_N5494_io_in_lo = {IN_CHANY_N27201_25,IN_CHANY_N27200_24,IN_CHANY_N27137_23,IN_CHANY_N27136_22,
    _CBMux_IPIN3_N5493_io_in_WIRE_1,IN_CHANY_N27118_4}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN4_N5494_io_in_hi = {IN_CHANY_N27237_79,IN_CHANY_N27236_78,IN_CHANY_N27227_43,IN_CHANY_N27226_42,
    IN_CHANY_N27203_33,IN_CHANY_N27202_32}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN5_N5495_io_in_lo = {IN_CHANY_N27200_24,IN_CHANY_N27137_23,IN_CHANY_N27136_22,IN_CHANY_N27129_15,
    IN_CHANY_N27128_14}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN5_N5495_io_in_hi = {_CBMux_IPIN1_N5491_io_in_WIRE_7,IN_CHANY_N27214_76,IN_CHANY_N27203_33,
    IN_CHANY_N27202_32,IN_CHANY_N27201_25}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN6_N5496_io_in_lo = {IN_CHANY_N27198_16,IN_CHANY_N27197_9,IN_CHANY_N27196_8,IN_CHANY_N27121_7,
    IN_CHANY_N27120_6}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN6_N5496_io_in_hi = {IN_CHANY_N27223_27,IN_CHANY_N27222_26,_CBMux_IPIN1_N5491_io_in_WIRE_7,
    IN_CHANY_N27214_76,IN_CHANY_N27199_17}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN7_N5497_io_in_lo = {IN_CHANY_N27219_11,IN_CHANY_N27218_10,IN_CHANY_N27195_1,IN_CHANY_N27194_0,
    _CBMux_IPIN1_N5491_io_in_WIRE_1,IN_CHANY_N27142_28}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN7_N5497_io_in_hi = {IN_CHANY_N27237_79,IN_CHANY_N27236_78,IN_CHANY_N27233_67,IN_CHANY_N27232_66,
    IN_CHANY_N27221_19,IN_CHANY_N27220_18}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN8_N5498_io_in_lo = {IN_CHANY_N27224_34,IN_CHANY_N27217_3,IN_CHANY_N27216_2,
    _CBMux_IPIN2_N5492_io_in_WIRE_1,IN_CHANY_N27134_20,_CBMux_IPIN3_N5493_io_in_WIRE_3,IN_CHANY_N27126_12}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN8_N5498_io_in_hi = {IN_CHANY_N27237_79,IN_CHANY_N27236_78,IN_CHANY_N27231_59,IN_CHANY_N27230_58,
    IN_CHANY_N27229_51,IN_CHANY_N27228_50,IN_CHANY_N27225_35}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN9_N5499_io_in_lo = {IN_CHANY_N27214_76,_CBMux_IPIN3_N5493_io_in_WIRE_7,IN_CHANY_N27150_36,
    IN_CHANY_N27145_31,IN_CHANY_N27144_30,_CBMux_IPIN3_N5493_io_in_WIRE_3,IN_CHANY_N27126_12}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN9_N5499_io_in_hi = {IN_CHANY_N27235_75,IN_CHANY_N27234_74,IN_CHANY_N27229_51,IN_CHANY_N27228_50,
    IN_CHANY_N27217_3,IN_CHANY_N27216_2,_CBMux_IPIN1_N5491_io_in_WIRE_7}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN10_N5500_io_in_lo = {IN_CHANY_N27150_36,IN_CHANY_N27145_31,IN_CHANY_N27144_30,IN_CHANY_N27137_23,
    IN_CHANY_N27136_22,_CBMux_IPIN3_N5493_io_in_WIRE_1,IN_CHANY_N27118_4}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN10_N5500_io_in_hi = {IN_CHANY_N27235_75,IN_CHANY_N27234_74,IN_CHANY_N27227_43,IN_CHANY_N27226_42,
    _CBMux_IPIN1_N5491_io_in_WIRE_7,IN_CHANY_N27214_76,_CBMux_IPIN3_N5493_io_in_WIRE_7}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN11_N5501_io_in_lo = {IN_CHANY_N27200_24,IN_CHANY_N27199_17,IN_CHANY_N27198_16,IN_CHANY_N27129_15,
    IN_CHANY_N27128_14}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN11_N5501_io_in_hi = {IN_CHANY_N27237_79,IN_CHANY_N27236_78,IN_CHANY_N27203_33,IN_CHANY_N27202_32,
    IN_CHANY_N27201_25}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN12_N5502_io_in_lo = {IN_CHANY_N27220_18,IN_CHANY_N27197_9,IN_CHANY_N27196_8,IN_CHANY_N27121_7,
    IN_CHANY_N27120_6}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN12_N5502_io_in_hi = {IN_CHANY_N27237_79,IN_CHANY_N27236_78,IN_CHANY_N27223_27,IN_CHANY_N27222_26,
    IN_CHANY_N27221_19}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN13_N5503_io_in_lo = {IN_CHANY_N27214_76,IN_CHANY_N27195_1,IN_CHANY_N27194_0,
    _CBMux_IPIN1_N5491_io_in_WIRE_1,IN_CHANY_N27142_28,_CBMux_IPIN2_N5492_io_in_WIRE_1,IN_CHANY_N27134_20}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN13_N5503_io_in_hi = {IN_CHANY_N27233_67,IN_CHANY_N27232_66,IN_CHANY_N27231_59,IN_CHANY_N27230_58,
    IN_CHANY_N27219_11,IN_CHANY_N27218_10,_CBMux_IPIN1_N5491_io_in_WIRE_7}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN14_N5504_io_in_lo = {_CBMux_IPIN1_N5491_io_in_WIRE_7,IN_CHANY_N27214_76,IN_CHANY_N27195_1,
    IN_CHANY_N27194_0,_CBMux_IPIN2_N5492_io_in_WIRE_1,IN_CHANY_N27134_20}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN15_N5505_io_in_lo = {IN_CHANY_N27217_3,IN_CHANY_N27216_2,IN_CHANY_N27145_31,IN_CHANY_N27144_30,
    _CBMux_IPIN3_N5493_io_in_WIRE_3,IN_CHANY_N27126_12}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN15_N5505_io_in_hi = {IN_CHANY_N27237_79,IN_CHANY_N27236_78,IN_CHANY_N27229_51,IN_CHANY_N27228_50,
    IN_CHANY_N27225_35,IN_CHANY_N27224_34}; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN16_N5506_io_in_lo = {IN_CHANX_N24003_15,IN_CHANX_N24002_14,IN_CHANX_N23995_7,IN_CHANX_N23994_6}; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN16_N5506_io_in_hi = {IN_CHANX_N24097_27,IN_CHANX_N24096_26,IN_CHANX_N24073_17,IN_CHANX_N24072_16}
    ; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN17_N5507_io_in_WIRE_1 = SBMux_C29_N24017_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire [4:0] CBMux_IPIN17_N5507_io_in_lo = {IN_CHANX_N24070_8,IN_CHANX_N24069_1,IN_CHANX_N24068_0,
    _CBMux_IPIN17_N5507_io_in_WIRE_1,IN_CHANX_N24016_28}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN17_N5507_io_in_hi = {IN_CHANX_N24107_67,IN_CHANX_N24106_66,IN_CHANX_N24095_19,IN_CHANX_N24094_18,
    IN_CHANX_N24071_9}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN18_N5508_io_in_WIRE_1 = SBMux_C21_N24009_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire [4:0] CBMux_IPIN18_N5508_io_in_lo = {IN_CHANX_N24092_10,IN_CHANX_N24091_3,IN_CHANX_N24090_2,
    _CBMux_IPIN18_N5508_io_in_WIRE_1,IN_CHANX_N24008_20}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN18_N5508_io_in_hi = {IN_CHANX_N24105_59,IN_CHANX_N24104_58,IN_CHANX_N24099_35,IN_CHANX_N24098_34,
    IN_CHANX_N24093_11}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN19_N5509_io_in_WIRE_1 = SBMux_C5_N23993_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN19_N5509_io_in_WIRE_3 = SBMux_C13_N24001_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire [6:0] CBMux_IPIN19_N5509_io_in_lo = {IN_CHANX_N24024_36,IN_CHANX_N24019_31,IN_CHANX_N24018_30,
    _CBMux_IPIN19_N5509_io_in_WIRE_3,IN_CHANX_N24000_12,_CBMux_IPIN19_N5509_io_in_WIRE_1,IN_CHANX_N23992_4}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN19_N5509_io_in_WIRE_7 = SBMux_C37_N24025_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire [6:0] CBMux_IPIN19_N5509_io_in_hi = {IN_CHANX_N24109_75,IN_CHANX_N24108_74,IN_CHANX_N24103_51,IN_CHANX_N24102_50,
    IN_CHANX_N24101_43,IN_CHANX_N24100_42,_CBMux_IPIN19_N5509_io_in_WIRE_7}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN20_N5510_io_in_lo = {IN_CHANX_N24074_24,IN_CHANX_N24011_23,IN_CHANX_N24010_22,
    _CBMux_IPIN19_N5509_io_in_WIRE_1,IN_CHANX_N23992_4}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN20_N5510_io_in_hi = {IN_CHANX_N24101_43,IN_CHANX_N24100_42,IN_CHANX_N24077_33,IN_CHANX_N24076_32,
    IN_CHANX_N24075_25}; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN21_N5511_io_in_lo = {IN_CHANX_N24011_23,IN_CHANX_N24010_22,IN_CHANX_N24003_15,IN_CHANX_N24002_14}
    ; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN21_N5511_io_in_hi = {IN_CHANX_N24077_33,IN_CHANX_N24076_32,IN_CHANX_N24075_25,IN_CHANX_N24074_24}
    ; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN22_N5512_io_in_lo = {IN_CHANX_N24071_9,IN_CHANX_N24070_8,IN_CHANX_N23995_7,IN_CHANX_N23994_6}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN23_N5513_io_in_lo = {IN_CHANX_N24092_10,IN_CHANX_N24069_1,IN_CHANX_N24068_0,
    _CBMux_IPIN17_N5507_io_in_WIRE_1,IN_CHANX_N24016_28}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN23_N5513_io_in_hi = {IN_CHANX_N24107_67,IN_CHANX_N24106_66,IN_CHANX_N24095_19,IN_CHANX_N24094_18,
    IN_CHANX_N24093_11}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN24_N5514_io_in_lo = {IN_CHANX_N24091_3,IN_CHANX_N24090_2,_CBMux_IPIN18_N5508_io_in_WIRE_1,
    IN_CHANX_N24008_20,_CBMux_IPIN19_N5509_io_in_WIRE_3,IN_CHANX_N24000_12}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN24_N5514_io_in_hi = {IN_CHANX_N24105_59,IN_CHANX_N24104_58,IN_CHANX_N24103_51,IN_CHANX_N24102_50,
    IN_CHANX_N24099_35,IN_CHANX_N24098_34}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN25_N5515_io_in_lo = {_CBMux_IPIN19_N5509_io_in_WIRE_7,IN_CHANX_N24024_36,IN_CHANX_N24019_31,
    IN_CHANX_N24018_30,_CBMux_IPIN19_N5509_io_in_WIRE_3,IN_CHANX_N24000_12}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN25_N5515_io_in_hi = {IN_CHANX_N24109_75,IN_CHANX_N24108_74,IN_CHANX_N24103_51,IN_CHANX_N24102_50,
    IN_CHANX_N24091_3,IN_CHANX_N24090_2}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN26_N5516_io_in_lo = {IN_CHANX_N24019_31,IN_CHANX_N24018_30,IN_CHANX_N24011_23,IN_CHANX_N24010_22,
    _CBMux_IPIN19_N5509_io_in_WIRE_1,IN_CHANX_N23992_4}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN26_N5516_io_in_hi = {IN_CHANX_N24109_75,IN_CHANX_N24108_74,IN_CHANX_N24101_43,IN_CHANX_N24100_42,
    _CBMux_IPIN19_N5509_io_in_WIRE_7,IN_CHANX_N24024_36}; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN27_N5517_io_in_lo = {IN_CHANX_N24073_17,IN_CHANX_N24072_16,IN_CHANX_N24003_15,IN_CHANX_N24002_14}
    ; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN28_N5518_io_in_hi = {IN_CHANX_N24097_27,IN_CHANX_N24096_26,IN_CHANX_N24095_19,IN_CHANX_N24094_18}
    ; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN29_N5519_io_in_lo = {IN_CHANX_N24069_1,IN_CHANX_N24068_0,_CBMux_IPIN17_N5507_io_in_WIRE_1,
    IN_CHANX_N24016_28,_CBMux_IPIN18_N5508_io_in_WIRE_1,IN_CHANX_N24008_20}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN29_N5519_io_in_hi = {IN_CHANX_N24107_67,IN_CHANX_N24106_66,IN_CHANX_N24105_59,IN_CHANX_N24104_58,
    IN_CHANX_N24093_11,IN_CHANX_N24092_10}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN30_N5520_io_in_lo = {IN_CHANX_N24092_10,IN_CHANX_N24069_1,IN_CHANX_N24068_0,
    _CBMux_IPIN18_N5508_io_in_WIRE_1,IN_CHANX_N24008_20}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN31_N5521_io_in_lo = {IN_CHANX_N24090_2,IN_CHANX_N24019_31,IN_CHANX_N24018_30,
    _CBMux_IPIN19_N5509_io_in_WIRE_3,IN_CHANX_N24000_12}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN31_N5521_io_in_hi = {IN_CHANX_N24103_51,IN_CHANX_N24102_50,IN_CHANX_N24099_35,IN_CHANX_N24098_34,
    IN_CHANX_N24091_3}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN32_N5522_io_in_lo = {IN_CHANX_N24024_36,IN_CHANX_N24011_23,IN_CHANX_N24010_22,
    _CBMux_IPIN19_N5509_io_in_WIRE_1,IN_CHANX_N23992_4}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN32_N5522_io_in_hi = {IN_CHANX_N24101_43,IN_CHANX_N24100_42,IN_CHANX_N24075_25,IN_CHANX_N24074_24,
    _CBMux_IPIN19_N5509_io_in_WIRE_7}; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN33_N5523_io_in_hi = {IN_CHANX_N24097_27,IN_CHANX_N24096_26,IN_CHANX_N24077_33,IN_CHANX_N24076_32}
    ; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN34_N5524_io_in_lo = {_CBMux_IPIN17_N5507_io_in_WIRE_1,IN_CHANX_N24016_28,IN_CHANX_N23995_7,
    IN_CHANX_N23994_6}; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN34_N5524_io_in_hi = {IN_CHANX_N24095_19,IN_CHANX_N24094_18,IN_CHANX_N24071_9,IN_CHANX_N24070_8}; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN36_N5526_io_in_lo = {IN_CHANX_N24069_1,IN_CHANX_N24068_0,_CBMux_IPIN18_N5508_io_in_WIRE_1,
    IN_CHANX_N24008_20}; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN36_N5526_io_in_hi = {IN_CHANX_N24099_35,IN_CHANX_N24098_34,IN_CHANX_N24093_11,IN_CHANX_N24092_10}
    ; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN37_N5527_io_in_lo = {IN_CHANX_N24024_36,IN_CHANX_N24019_31,IN_CHANX_N24018_30,
    _CBMux_IPIN19_N5509_io_in_WIRE_3,IN_CHANX_N24000_12}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN37_N5527_io_in_hi = {IN_CHANX_N24103_51,IN_CHANX_N24102_50,IN_CHANX_N24091_3,IN_CHANX_N24090_2,
    _CBMux_IPIN19_N5509_io_in_WIRE_7}; // @[TileFull.scala 166:8]
  wire  _SBMux_C5_N23993_O_3_C_6_io_in_WIRE_1 = logicBlock_OPIN_83; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C5_N23993_O_3_C_6_io_in_WIRE_0 = logicBlock_OPIN_81; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C5_N23993_O_3_C_6_io_in_WIRE_2 = logicBlock_OPIN_86; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C5_N23993_O_3_C_6_io_in_lo = {IN_CHANX_N24113_5,_SBMux_C5_N23993_O_3_C_6_io_in_WIRE_2,
    _SBMux_C5_N23993_O_3_C_6_io_in_WIRE_1,_SBMux_C5_N23993_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C5_N23993_O_3_C_6_io_in_hi = {IN_CHANY_N27239_5,IN_CHANY_N27223_27,IN_CHANY_N27214_76,
    IN_CHANY_N27200_24,IN_CHANY_N27195_1}; // @[TileFull.scala 183:11]
  wire  _SBMux_C13_N24001_O_3_C_6_io_in_WIRE_1 = logicBlock_OPIN_84; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C13_N24001_O_3_C_6_io_in_lo = {IN_CHANX_N24115_13,_SBMux_C5_N23993_O_3_C_6_io_in_WIRE_2,
    _SBMux_C13_N24001_O_3_C_6_io_in_WIRE_1,_SBMux_C5_N23993_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C13_N24001_O_3_C_6_io_in_hi = {IN_CHANY_N27257_77,IN_CHANY_N27222_26,IN_CHANY_N27201_25,
    IN_CHANY_N27194_0,IN_CHANY_N27118_4}; // @[TileFull.scala 183:11]
  wire  _SBMux_C21_N24009_O_3_C_6_io_in_WIRE_0 = logicBlock_OPIN_82; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C21_N24009_O_3_C_6_io_in_WIRE_2 = logicBlock_OPIN_87; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C21_N24009_O_3_C_6_io_in_lo = {IN_CHANX_N24117_21,_SBMux_C21_N24009_O_3_C_6_io_in_WIRE_2,
    _SBMux_C13_N24001_O_3_C_6_io_in_WIRE_1,_SBMux_C21_N24009_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C21_N24009_O_3_C_6_io_in_hi = {IN_CHANY_N27255_69,IN_CHANY_N27216_2,IN_CHANY_N27144_30,
    IN_CHANY_N27137_23,IN_CHANY_N27126_12}; // @[TileFull.scala 183:11]
  wire  _SBMux_C29_N24017_O_3_C_6_io_in_WIRE_1 = logicBlock_OPIN_85; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C29_N24017_O_3_C_6_io_in_lo = {IN_CHANX_N24119_29,_SBMux_C21_N24009_O_3_C_6_io_in_WIRE_2,
    _SBMux_C29_N24017_O_3_C_6_io_in_WIRE_1,_SBMux_C21_N24009_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C29_N24017_O_3_C_6_io_in_hi = {IN_CHANY_N27253_61,IN_CHANY_N27221_19,IN_CHANY_N27202_32,
    IN_CHANY_N27134_20,IN_CHANY_N27120_6}; // @[TileFull.scala 183:11]
  wire  _SBMux_C37_N24025_O_3_C_6_io_in_WIRE_2 = logicBlock_OPIN_88; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C37_N24025_O_3_C_6_io_in_lo = {IN_CHANX_N24121_37,_SBMux_C37_N24025_O_3_C_6_io_in_WIRE_2,
    _SBMux_C29_N24017_O_3_C_6_io_in_WIRE_1,_SBMux_C5_N23993_O_3_C_6_io_in_WIRE_1}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C37_N24025_O_3_C_6_io_in_hi = {IN_CHANY_N27251_53,IN_CHANY_N27224_34,IN_CHANY_N27199_17,
    IN_CHANY_N27196_8,IN_CHANY_N27142_28}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C45_N24033_O_4_C_5_io_in_lo = {_SBMux_C21_N24009_O_3_C_6_io_in_WIRE_2,
    _SBMux_C29_N24017_O_3_C_6_io_in_WIRE_1,_SBMux_C5_N23993_O_3_C_6_io_in_WIRE_1,_SBMux_C5_N23993_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C45_N24033_O_4_C_5_io_in_hi = {IN_CHANY_N27249_45,IN_CHANY_N27218_10,IN_CHANY_N27150_36,
    IN_CHANY_N27129_15,IN_CHANX_N24123_45}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C53_N24041_O_4_C_5_io_in_hi = {IN_CHANY_N27247_37,IN_CHANY_N27219_11,IN_CHANY_N27158_44,
    IN_CHANY_N27128_14,IN_CHANX_N24125_53}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C61_N24049_O_4_C_6_io_in_lo = {IN_CHANX_N24127_61,_SBMux_C37_N24025_O_3_C_6_io_in_WIRE_2,
    _SBMux_C5_N23993_O_3_C_6_io_in_WIRE_2,_SBMux_C13_N24001_O_3_C_6_io_in_WIRE_1,_SBMux_C21_N24009_O_3_C_6_io_in_WIRE_0}
    ; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C61_N24049_O_4_C_6_io_in_hi = {IN_CHANY_N27245_29,IN_CHANY_N27225_35,IN_CHANY_N27198_16,
    IN_CHANY_N27197_9,IN_CHANY_N27166_52}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C69_N24057_O_3_C_6_io_in_lo = {IN_CHANX_N24129_69,_SBMux_C5_N23993_O_3_C_6_io_in_WIRE_2,
    _SBMux_C13_N24001_O_3_C_6_io_in_WIRE_1,_SBMux_C21_N24009_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C69_N24057_O_3_C_6_io_in_hi = {IN_CHANY_N27243_21,IN_CHANY_N27220_18,IN_CHANY_N27203_33,
    IN_CHANY_N27174_60,IN_CHANY_N27121_7}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C77_N24089_O_0_C_6_io_in_lo = {IN_CHANY_N27145_31,IN_CHANY_N27136_22,IN_CHANX_N24131_77}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C77_N24089_O_0_C_6_io_in_hi = {IN_CHANY_N27241_13,IN_CHANY_N27217_3,IN_CHANY_N27182_68}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C4_N24112_O_3_C_5_io_in_lo = {IN_CHANX_N23992_4,IN_OPIN_N8016_86,IN_OPIN_N8013_83,IN_OPIN_N8011_81}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C4_N24112_O_3_C_5_io_in_hi = {IN_CHANY_N27257_77,IN_CHANY_N27201_25,IN_CHANY_N27182_68,
    IN_CHANY_N27136_22}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C12_N24114_O_3_C_6_io_in_lo = {IN_CHANX_N24000_12,IN_OPIN_N8016_86,IN_OPIN_N8014_84,IN_OPIN_N8011_81}
    ; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C12_N24114_O_3_C_6_io_in_hi = {IN_CHANY_N27239_5,IN_CHANY_N27223_27,IN_CHANY_N27220_18,
    IN_CHANY_N27195_1,IN_CHANY_N27174_60}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C20_N24116_O_3_C_6_io_in_lo = {IN_CHANX_N24008_20,IN_OPIN_N8017_87,IN_OPIN_N8014_84,IN_OPIN_N8012_82}
    ; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C20_N24116_O_3_C_6_io_in_hi = {IN_CHANY_N27241_13,IN_CHANY_N27217_3,IN_CHANY_N27198_16,
    IN_CHANY_N27166_52,IN_CHANY_N27145_31}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C28_N24118_O_3_C_6_io_in_lo = {IN_CHANX_N24016_28,IN_OPIN_N8017_87,IN_OPIN_N8015_85,IN_OPIN_N8012_82}
    ; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C28_N24118_O_3_C_6_io_in_hi = {IN_CHANY_N27243_21,IN_CHANY_N27203_33,IN_CHANY_N27158_44,
    IN_CHANY_N27128_14,IN_CHANY_N27121_7}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C36_N24120_O_3_C_6_io_in_lo = {IN_CHANX_N24024_36,IN_OPIN_N8018_88,IN_OPIN_N8015_85,IN_OPIN_N8013_83}
    ; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C36_N24120_O_3_C_6_io_in_hi = {IN_CHANY_N27245_29,IN_CHANY_N27225_35,IN_CHANY_N27218_10,
    IN_CHANY_N27197_9,IN_CHANY_N27150_36}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C44_N24122_O_4_C_5_io_in_lo = {IN_OPIN_N8017_87,IN_OPIN_N8015_85,IN_OPIN_N8013_83,IN_OPIN_N8011_81}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C44_N24122_O_4_C_5_io_in_hi = {IN_CHANY_N27247_37,IN_CHANY_N27219_11,IN_CHANY_N27196_8,
    IN_CHANY_N27142_28,IN_CHANX_N24032_44}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C52_N24124_O_4_C_5_io_in_hi = {IN_CHANY_N27249_45,IN_CHANY_N27134_20,IN_CHANY_N27129_15,
    IN_CHANY_N27120_6,IN_CHANX_N24040_52}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C60_N24126_O_4_C_5_io_in_lo = {IN_OPIN_N8018_88,IN_OPIN_N8016_86,IN_OPIN_N8014_84,IN_OPIN_N8012_82}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C60_N24126_O_4_C_5_io_in_hi = {IN_CHANY_N27251_53,IN_CHANY_N27216_2,IN_CHANY_N27199_17,
    IN_CHANY_N27126_12,IN_CHANX_N24048_60}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C68_N24128_O_3_C_5_io_in_lo = {IN_CHANX_N24056_68,IN_OPIN_N8016_86,IN_OPIN_N8014_84,IN_OPIN_N8012_82}
    ; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C68_N24128_O_3_C_5_io_in_hi = {IN_CHANY_N27253_61,IN_CHANY_N27221_19,IN_CHANY_N27194_0,
    IN_CHANY_N27118_4}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C76_N24130_O_0_C_4_io_in_lo = {IN_CHANY_N27137_23,IN_CHANX_N24088_76}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C76_N24130_O_0_C_4_io_in_hi = {IN_CHANY_N27255_69,IN_CHANY_N27214_76}; // @[TileFull.scala 183:11]
  wire  _SBMux_C5_N27119_O_4_C_6_io_in_WIRE_1 = logicBlock_OPIN_75; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C5_N27119_O_4_C_6_io_in_WIRE_0 = logicBlock_OPIN_73; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C5_N27119_O_4_C_6_io_in_WIRE_3 = logicBlock_OPIN_80; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C5_N27119_O_4_C_6_io_in_WIRE_2 = logicBlock_OPIN_78; // @[TileFull.scala 174:{37,37}]
  wire [4:0] SBMux_C5_N27119_O_4_C_6_io_in_lo = {IN_CHANX_N24000_12,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_3,
    _SBMux_C5_N27119_O_4_C_6_io_in_WIRE_2,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_1,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C5_N27119_O_4_C_6_io_in_hi = {IN_CHANY_N27239_5,IN_CHANX_N24129_69,IN_CHANX_N24090_2,
    IN_CHANX_N24018_30,IN_CHANX_N24011_23}; // @[TileFull.scala 183:11]
  wire  _SBMux_C13_N27127_O_3_C_6_io_in_WIRE_1 = logicBlock_OPIN_76; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C13_N27127_O_3_C_6_io_in_lo = {IN_CHANX_N23994_6,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_2,
    _SBMux_C13_N27127_O_3_C_6_io_in_WIRE_1,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C13_N27127_O_3_C_6_io_in_hi = {IN_CHANY_N27241_13,IN_CHANX_N24127_61,IN_CHANX_N24095_19,
    IN_CHANX_N24076_32,IN_CHANX_N24008_20}; // @[TileFull.scala 183:11]
  wire  _SBMux_C21_N27135_O_3_C_6_io_in_WIRE_0 = logicBlock_OPIN_74; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C21_N27135_O_3_C_6_io_in_WIRE_2 = logicBlock_OPIN_79; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C21_N27135_O_3_C_6_io_in_lo = {IN_CHANX_N24016_28,_SBMux_C21_N27135_O_3_C_6_io_in_WIRE_2,
    _SBMux_C13_N27127_O_3_C_6_io_in_WIRE_1,_SBMux_C21_N27135_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C21_N27135_O_3_C_6_io_in_hi = {IN_CHANY_N27243_21,IN_CHANX_N24125_53,IN_CHANX_N24098_34,
    IN_CHANX_N24073_17,IN_CHANX_N24070_8}; // @[TileFull.scala 183:11]
  wire  _SBMux_C29_N27143_O_3_C_5_io_in_WIRE_1 = logicBlock_OPIN_77; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C29_N27143_O_3_C_5_io_in_lo = {IN_CHANX_N24003_15,_SBMux_C21_N27135_O_3_C_6_io_in_WIRE_2,
    _SBMux_C29_N27143_O_3_C_5_io_in_WIRE_1,_SBMux_C21_N27135_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C29_N27143_O_3_C_5_io_in_hi = {IN_CHANY_N27245_29,IN_CHANX_N24123_45,IN_CHANX_N24092_10,
    IN_CHANX_N24024_36}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C37_N27151_O_3_C_5_io_in_lo = {IN_CHANX_N24002_14,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_3,
    _SBMux_C29_N27143_O_3_C_5_io_in_WIRE_1,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_1}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C37_N27151_O_3_C_5_io_in_hi = {IN_CHANY_N27247_37,IN_CHANX_N24121_37,IN_CHANX_N24093_11,
    IN_CHANX_N24032_44}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C45_N27159_O_4_C_5_io_in_lo = {_SBMux_C21_N27135_O_3_C_6_io_in_WIRE_2,
    _SBMux_C29_N27143_O_3_C_5_io_in_WIRE_1,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_1,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C45_N27159_O_4_C_5_io_in_hi = {IN_CHANY_N27249_45,IN_CHANX_N24119_29,IN_CHANX_N24072_16,
    IN_CHANX_N24071_9,IN_CHANX_N24040_52}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C53_N27167_O_4_C_5_io_in_hi = {IN_CHANY_N27251_53,IN_CHANX_N24117_21,IN_CHANX_N24094_18,
    IN_CHANX_N24048_60,IN_CHANX_N23995_7}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C61_N27175_O_4_C_5_io_in_lo = {_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_3,
    _SBMux_C5_N27119_O_4_C_6_io_in_WIRE_2,_SBMux_C13_N27127_O_3_C_6_io_in_WIRE_1,_SBMux_C21_N27135_O_3_C_6_io_in_WIRE_0}
    ; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C61_N27175_O_4_C_5_io_in_hi = {IN_CHANY_N27253_61,IN_CHANX_N24115_13,IN_CHANX_N24091_3,
    IN_CHANX_N24056_68,IN_CHANX_N24010_22}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C69_N27183_O_4_C_5_io_in_hi = {IN_CHANY_N27255_69,IN_CHANX_N24113_5,IN_CHANX_N24088_76,
    IN_CHANX_N24074_24,IN_CHANX_N24069_1}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C77_N27215_O_3_C_5_io_in_lo = {IN_CHANX_N23992_4,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_1,
    _SBMux_C21_N27135_O_3_C_6_io_in_WIRE_0,_SBMux_C5_N27119_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C77_N27215_O_3_C_5_io_in_hi = {IN_CHANY_N27257_77,IN_CHANX_N24131_77,IN_CHANX_N24096_26,
    IN_CHANX_N24068_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C4_N27238_O_4_C_7_io_in_lo = {IN_CHANX_N23992_4,IN_OPIN_N5814_80,IN_OPIN_N5812_78,IN_OPIN_N5809_75,
    IN_OPIN_N5807_73}; // @[TileFull.scala 183:11]
  wire [5:0] SBMux_C4_N27238_O_4_C_7_io_in_hi = {IN_CHANY_N27118_4,IN_CHANX_N24115_13,IN_CHANX_N24096_26,
    IN_CHANX_N24091_3,IN_CHANX_N24068_0,IN_CHANX_N24019_31}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C12_N27240_O_3_C_6_io_in_lo = {IN_CHANX_N23995_7,IN_OPIN_N5812_78,IN_OPIN_N5810_76,IN_OPIN_N5807_73}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C12_N27240_O_3_C_6_io_in_hi = {IN_CHANY_N27126_12,IN_CHANX_N24117_21,IN_CHANX_N24088_76,
    IN_CHANX_N24077_33,IN_CHANX_N24074_24}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C20_N27242_O_3_C_6_io_in_lo = {IN_CHANX_N24010_22,IN_OPIN_N5813_79,IN_OPIN_N5810_76,IN_OPIN_N5808_74}
    ; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C20_N27242_O_3_C_6_io_in_hi = {IN_CHANY_N27134_20,IN_CHANX_N24119_29,IN_CHANX_N24099_35,
    IN_CHANX_N24071_9,IN_CHANX_N24056_68}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C28_N27244_O_3_C_5_io_in_lo = {IN_CHANX_N24048_60,IN_OPIN_N5813_79,IN_OPIN_N5811_77,IN_OPIN_N5808_74}
    ; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C28_N27244_O_3_C_5_io_in_hi = {IN_CHANY_N27142_28,IN_CHANX_N24121_37,IN_CHANX_N24094_18,
    IN_CHANX_N24093_11}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C36_N27246_O_3_C_5_io_in_lo = {IN_CHANX_N24003_15,IN_OPIN_N5814_80,IN_OPIN_N5811_77,IN_OPIN_N5809_75}
    ; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C36_N27246_O_3_C_5_io_in_hi = {IN_CHANY_N27150_36,IN_CHANX_N24123_45,IN_CHANX_N24072_16,
    IN_CHANX_N24040_52}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C44_N27248_O_4_C_5_io_in_lo = {IN_OPIN_N5813_79,IN_OPIN_N5811_77,IN_OPIN_N5809_75,IN_OPIN_N5807_73}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C44_N27248_O_4_C_5_io_in_hi = {IN_CHANY_N27158_44,IN_CHANX_N24125_53,IN_CHANX_N24073_17,
    IN_CHANX_N24032_44,IN_CHANX_N24002_14}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C52_N27250_O_4_C_5_io_in_hi = {IN_CHANY_N27166_52,IN_CHANX_N24127_61,IN_CHANX_N24095_19,
    IN_CHANX_N24092_10,IN_CHANX_N24024_36}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C60_N27252_O_4_C_6_io_in_lo = {IN_CHANX_N24011_23,IN_OPIN_N5814_80,IN_OPIN_N5812_78,IN_OPIN_N5810_76,
    IN_OPIN_N5808_74}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C60_N27252_O_4_C_6_io_in_hi = {IN_CHANY_N27174_60,IN_CHANX_N24129_69,IN_CHANX_N24098_34,
    IN_CHANX_N24070_8,IN_CHANX_N24016_28}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C68_N27254_O_4_C_6_io_in_lo = {IN_CHANX_N23994_6,IN_OPIN_N5814_80,IN_OPIN_N5812_78,IN_OPIN_N5810_76,
    IN_OPIN_N5808_74}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C68_N27254_O_4_C_6_io_in_hi = {IN_CHANY_N27182_68,IN_CHANX_N24131_77,IN_CHANX_N24076_32,
    IN_CHANX_N24075_25,IN_CHANX_N24008_20}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C76_N27256_O_3_C_7_io_in_lo = {IN_CHANX_N24018_30,IN_CHANX_N24000_12,IN_OPIN_N5809_75,
    IN_OPIN_N5808_74,IN_OPIN_N5807_73}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C76_N27256_O_3_C_7_io_in_hi = {IN_CHANY_N27214_76,IN_CHANX_N24113_5,IN_CHANX_N24097_27,
    IN_CHANX_N24090_2,IN_CHANX_N24069_1}; // @[TileFull.scala 183:11]
  CLBlut4N10Alu logicBlock ( // @[TileFull.scala 47:37]
    .IPIN_0(logicBlock_IPIN_0),
    .IPIN_1(logicBlock_IPIN_1),
    .IPIN_2(logicBlock_IPIN_2),
    .IPIN_3(logicBlock_IPIN_3),
    .IPIN_4(logicBlock_IPIN_4),
    .IPIN_5(logicBlock_IPIN_5),
    .IPIN_6(logicBlock_IPIN_6),
    .IPIN_7(logicBlock_IPIN_7),
    .IPIN_8(logicBlock_IPIN_8),
    .IPIN_9(logicBlock_IPIN_9),
    .IPIN_10(logicBlock_IPIN_10),
    .IPIN_11(logicBlock_IPIN_11),
    .IPIN_12(logicBlock_IPIN_12),
    .IPIN_13(logicBlock_IPIN_13),
    .IPIN_14(logicBlock_IPIN_14),
    .IPIN_15(logicBlock_IPIN_15),
    .IPIN_16(logicBlock_IPIN_16),
    .IPIN_17(logicBlock_IPIN_17),
    .IPIN_18(logicBlock_IPIN_18),
    .IPIN_19(logicBlock_IPIN_19),
    .IPIN_20(logicBlock_IPIN_20),
    .IPIN_21(logicBlock_IPIN_21),
    .IPIN_22(logicBlock_IPIN_22),
    .IPIN_23(logicBlock_IPIN_23),
    .IPIN_24(logicBlock_IPIN_24),
    .IPIN_25(logicBlock_IPIN_25),
    .IPIN_26(logicBlock_IPIN_26),
    .IPIN_27(logicBlock_IPIN_27),
    .IPIN_28(logicBlock_IPIN_28),
    .IPIN_29(logicBlock_IPIN_29),
    .IPIN_30(logicBlock_IPIN_30),
    .IPIN_31(logicBlock_IPIN_31),
    .IPIN_32(logicBlock_IPIN_32),
    .IPIN_33(logicBlock_IPIN_33),
    .IPIN_34(logicBlock_IPIN_34),
    .IPIN_35(logicBlock_IPIN_35),
    .IPIN_36(logicBlock_IPIN_36),
    .IPIN_37(logicBlock_IPIN_37),
    .IPIN_38(logicBlock_IPIN_38),
    .IPIN_39(logicBlock_IPIN_39),
    .IPIN_40(logicBlock_IPIN_40),
    .IPIN_41(logicBlock_IPIN_41),
    .IPIN_42(logicBlock_IPIN_42),
    .IPIN_43(logicBlock_IPIN_43),
    .IPIN_44(logicBlock_IPIN_44),
    .IPIN_45(logicBlock_IPIN_45),
    .IPIN_46(logicBlock_IPIN_46),
    .IPIN_47(logicBlock_IPIN_47),
    .IPIN_48(logicBlock_IPIN_48),
    .IPIN_49(logicBlock_IPIN_49),
    .IPIN_50(logicBlock_IPIN_50),
    .IPIN_51(logicBlock_IPIN_51),
    .IPIN_52(logicBlock_IPIN_52),
    .IPIN_53(logicBlock_IPIN_53),
    .IPIN_54(logicBlock_IPIN_54),
    .IPIN_55(logicBlock_IPIN_55),
    .IPIN_56(logicBlock_IPIN_56),
    .IPIN_57(logicBlock_IPIN_57),
    .IPIN_58(logicBlock_IPIN_58),
    .IPIN_59(logicBlock_IPIN_59),
    .IPIN_60(logicBlock_IPIN_60),
    .IPIN_61(logicBlock_IPIN_61),
    .IPIN_62(logicBlock_IPIN_62),
    .IPIN_63(logicBlock_IPIN_63),
    .IPIN_64(logicBlock_IPIN_64),
    .IPIN_65(logicBlock_IPIN_65),
    .IPIN_66(logicBlock_IPIN_66),
    .IPIN_67(logicBlock_IPIN_67),
    .IPIN_68(logicBlock_IPIN_68),
    .IPIN_69(logicBlock_IPIN_69),
    .IPIN_70(logicBlock_IPIN_70),
    .IPIN_71(logicBlock_IPIN_71),
    .OPIN_73(logicBlock_OPIN_73),
    .OPIN_74(logicBlock_OPIN_74),
    .OPIN_75(logicBlock_OPIN_75),
    .OPIN_76(logicBlock_OPIN_76),
    .OPIN_77(logicBlock_OPIN_77),
    .OPIN_78(logicBlock_OPIN_78),
    .OPIN_79(logicBlock_OPIN_79),
    .OPIN_80(logicBlock_OPIN_80),
    .OPIN_81(logicBlock_OPIN_81),
    .OPIN_82(logicBlock_OPIN_82),
    .OPIN_83(logicBlock_OPIN_83),
    .OPIN_84(logicBlock_OPIN_84),
    .OPIN_85(logicBlock_OPIN_85),
    .OPIN_86(logicBlock_OPIN_86),
    .OPIN_87(logicBlock_OPIN_87),
    .OPIN_88(logicBlock_OPIN_88),
    .OPIN_89(logicBlock_OPIN_89),
    .OPIN_90(logicBlock_OPIN_90),
    .OPIN_91(logicBlock_OPIN_91),
    .OPIN_92(logicBlock_OPIN_92),
    .OPIN_93(logicBlock_OPIN_93),
    .OPIN_94(logicBlock_OPIN_94),
    .OPIN_95(logicBlock_OPIN_95),
    .OPIN_96(logicBlock_OPIN_96),
    .OPIN_97(logicBlock_OPIN_97),
    .OPIN_98(logicBlock_OPIN_98),
    .OPIN_99(logicBlock_OPIN_99),
    .OPIN_100(logicBlock_OPIN_100),
    .OPIN_101(logicBlock_OPIN_101),
    .OPIN_102(logicBlock_OPIN_102),
    .OPIN_103(logicBlock_OPIN_103),
    .OPIN_104(logicBlock_OPIN_104),
    .OPIN_105(logicBlock_OPIN_105),
    .OPIN_106(logicBlock_OPIN_106),
    .OPIN_107(logicBlock_OPIN_107),
    .OPIN_108(logicBlock_OPIN_108),
    .OPIN_109(logicBlock_OPIN_109),
    .OPIN_110(logicBlock_OPIN_110),
    .OPIN_111(logicBlock_OPIN_111),
    .OPIN_112(logicBlock_OPIN_112),
    .OPIN_113(logicBlock_OPIN_113),
    .OPIN_114(logicBlock_OPIN_114),
    .OPIN_115(logicBlock_OPIN_115),
    .OPIN_116(logicBlock_OPIN_116),
    .OPIN_117(logicBlock_OPIN_117),
    .OPIN_118(logicBlock_OPIN_118),
    .OPIN_119(logicBlock_OPIN_119),
    .OPIN_120(logicBlock_OPIN_120),
    .clock(logicBlock_clock),
    .reset(logicBlock_reset),
    .configBits(logicBlock_configBits),
    .gndLBouts(logicBlock_gndLBouts)
  );
  ScanConf_Tile_3_3_clbalutile configBlock ( // @[TileFull.scala 61:31]
    .clock(configBlock_clock),
    .ioBundle_confOut(configBlock_ioBundle_confOut),
    .ioBundle_scan_in(configBlock_ioBundle_scan_in),
    .ioBundle_scan_en(configBlock_ioBundle_scan_en),
    .ioBundle_scan_out(configBlock_ioBundle_scan_out)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN0_N5490 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN0_N5490_io_in),
    .io_config(CBMux_IPIN0_N5490_io_config),
    .io_out(CBMux_IPIN0_N5490_io_out),
    .io_loopBreak(CBMux_IPIN0_N5490_io_loopBreak),
    .io_cnstClk(CBMux_IPIN0_N5490_io_cnstClk),
    .io_arst(CBMux_IPIN0_N5490_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN1_N5491 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN1_N5491_io_in),
    .io_config(CBMux_IPIN1_N5491_io_config),
    .io_out(CBMux_IPIN1_N5491_io_out),
    .io_loopBreak(CBMux_IPIN1_N5491_io_loopBreak),
    .io_cnstClk(CBMux_IPIN1_N5491_io_cnstClk),
    .io_arst(CBMux_IPIN1_N5491_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN2_N5492 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN2_N5492_io_in),
    .io_config(CBMux_IPIN2_N5492_io_config),
    .io_out(CBMux_IPIN2_N5492_io_out),
    .io_loopBreak(CBMux_IPIN2_N5492_io_loopBreak),
    .io_cnstClk(CBMux_IPIN2_N5492_io_cnstClk),
    .io_arst(CBMux_IPIN2_N5492_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN3_N5493 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN3_N5493_io_in),
    .io_config(CBMux_IPIN3_N5493_io_config),
    .io_out(CBMux_IPIN3_N5493_io_out),
    .io_loopBreak(CBMux_IPIN3_N5493_io_loopBreak),
    .io_cnstClk(CBMux_IPIN3_N5493_io_cnstClk),
    .io_arst(CBMux_IPIN3_N5493_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN4_N5494 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN4_N5494_io_in),
    .io_config(CBMux_IPIN4_N5494_io_config),
    .io_out(CBMux_IPIN4_N5494_io_out),
    .io_loopBreak(CBMux_IPIN4_N5494_io_loopBreak),
    .io_cnstClk(CBMux_IPIN4_N5494_io_cnstClk),
    .io_arst(CBMux_IPIN4_N5494_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN5_N5495 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN5_N5495_io_in),
    .io_config(CBMux_IPIN5_N5495_io_config),
    .io_out(CBMux_IPIN5_N5495_io_out),
    .io_loopBreak(CBMux_IPIN5_N5495_io_loopBreak),
    .io_cnstClk(CBMux_IPIN5_N5495_io_cnstClk),
    .io_arst(CBMux_IPIN5_N5495_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN6_N5496 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN6_N5496_io_in),
    .io_config(CBMux_IPIN6_N5496_io_config),
    .io_out(CBMux_IPIN6_N5496_io_out),
    .io_loopBreak(CBMux_IPIN6_N5496_io_loopBreak),
    .io_cnstClk(CBMux_IPIN6_N5496_io_cnstClk),
    .io_arst(CBMux_IPIN6_N5496_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN7_N5497 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN7_N5497_io_in),
    .io_config(CBMux_IPIN7_N5497_io_config),
    .io_out(CBMux_IPIN7_N5497_io_out),
    .io_loopBreak(CBMux_IPIN7_N5497_io_loopBreak),
    .io_cnstClk(CBMux_IPIN7_N5497_io_cnstClk),
    .io_arst(CBMux_IPIN7_N5497_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN8_N5498 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN8_N5498_io_in),
    .io_config(CBMux_IPIN8_N5498_io_config),
    .io_out(CBMux_IPIN8_N5498_io_out),
    .io_loopBreak(CBMux_IPIN8_N5498_io_loopBreak),
    .io_cnstClk(CBMux_IPIN8_N5498_io_cnstClk),
    .io_arst(CBMux_IPIN8_N5498_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN9_N5499 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN9_N5499_io_in),
    .io_config(CBMux_IPIN9_N5499_io_config),
    .io_out(CBMux_IPIN9_N5499_io_out),
    .io_loopBreak(CBMux_IPIN9_N5499_io_loopBreak),
    .io_cnstClk(CBMux_IPIN9_N5499_io_cnstClk),
    .io_arst(CBMux_IPIN9_N5499_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN10_N5500 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN10_N5500_io_in),
    .io_config(CBMux_IPIN10_N5500_io_config),
    .io_out(CBMux_IPIN10_N5500_io_out),
    .io_loopBreak(CBMux_IPIN10_N5500_io_loopBreak),
    .io_cnstClk(CBMux_IPIN10_N5500_io_cnstClk),
    .io_arst(CBMux_IPIN10_N5500_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN11_N5501 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN11_N5501_io_in),
    .io_config(CBMux_IPIN11_N5501_io_config),
    .io_out(CBMux_IPIN11_N5501_io_out),
    .io_loopBreak(CBMux_IPIN11_N5501_io_loopBreak),
    .io_cnstClk(CBMux_IPIN11_N5501_io_cnstClk),
    .io_arst(CBMux_IPIN11_N5501_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN12_N5502 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN12_N5502_io_in),
    .io_config(CBMux_IPIN12_N5502_io_config),
    .io_out(CBMux_IPIN12_N5502_io_out),
    .io_loopBreak(CBMux_IPIN12_N5502_io_loopBreak),
    .io_cnstClk(CBMux_IPIN12_N5502_io_cnstClk),
    .io_arst(CBMux_IPIN12_N5502_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN13_N5503 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN13_N5503_io_in),
    .io_config(CBMux_IPIN13_N5503_io_config),
    .io_out(CBMux_IPIN13_N5503_io_out),
    .io_loopBreak(CBMux_IPIN13_N5503_io_loopBreak),
    .io_cnstClk(CBMux_IPIN13_N5503_io_cnstClk),
    .io_arst(CBMux_IPIN13_N5503_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN14_N5504 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN14_N5504_io_in),
    .io_config(CBMux_IPIN14_N5504_io_config),
    .io_out(CBMux_IPIN14_N5504_io_out),
    .io_loopBreak(CBMux_IPIN14_N5504_io_loopBreak),
    .io_cnstClk(CBMux_IPIN14_N5504_io_cnstClk),
    .io_arst(CBMux_IPIN14_N5504_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN15_N5505 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN15_N5505_io_in),
    .io_config(CBMux_IPIN15_N5505_io_config),
    .io_out(CBMux_IPIN15_N5505_io_out),
    .io_loopBreak(CBMux_IPIN15_N5505_io_loopBreak),
    .io_cnstClk(CBMux_IPIN15_N5505_io_cnstClk),
    .io_arst(CBMux_IPIN15_N5505_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN16_N5506 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN16_N5506_io_in),
    .io_config(CBMux_IPIN16_N5506_io_config),
    .io_out(CBMux_IPIN16_N5506_io_out),
    .io_loopBreak(CBMux_IPIN16_N5506_io_loopBreak),
    .io_cnstClk(CBMux_IPIN16_N5506_io_cnstClk),
    .io_arst(CBMux_IPIN16_N5506_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN17_N5507 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN17_N5507_io_in),
    .io_config(CBMux_IPIN17_N5507_io_config),
    .io_out(CBMux_IPIN17_N5507_io_out),
    .io_loopBreak(CBMux_IPIN17_N5507_io_loopBreak),
    .io_cnstClk(CBMux_IPIN17_N5507_io_cnstClk),
    .io_arst(CBMux_IPIN17_N5507_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN18_N5508 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN18_N5508_io_in),
    .io_config(CBMux_IPIN18_N5508_io_config),
    .io_out(CBMux_IPIN18_N5508_io_out),
    .io_loopBreak(CBMux_IPIN18_N5508_io_loopBreak),
    .io_cnstClk(CBMux_IPIN18_N5508_io_cnstClk),
    .io_arst(CBMux_IPIN18_N5508_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN19_N5509 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN19_N5509_io_in),
    .io_config(CBMux_IPIN19_N5509_io_config),
    .io_out(CBMux_IPIN19_N5509_io_out),
    .io_loopBreak(CBMux_IPIN19_N5509_io_loopBreak),
    .io_cnstClk(CBMux_IPIN19_N5509_io_cnstClk),
    .io_arst(CBMux_IPIN19_N5509_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN20_N5510 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN20_N5510_io_in),
    .io_config(CBMux_IPIN20_N5510_io_config),
    .io_out(CBMux_IPIN20_N5510_io_out),
    .io_loopBreak(CBMux_IPIN20_N5510_io_loopBreak),
    .io_cnstClk(CBMux_IPIN20_N5510_io_cnstClk),
    .io_arst(CBMux_IPIN20_N5510_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN21_N5511 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN21_N5511_io_in),
    .io_config(CBMux_IPIN21_N5511_io_config),
    .io_out(CBMux_IPIN21_N5511_io_out),
    .io_loopBreak(CBMux_IPIN21_N5511_io_loopBreak),
    .io_cnstClk(CBMux_IPIN21_N5511_io_cnstClk),
    .io_arst(CBMux_IPIN21_N5511_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN22_N5512 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN22_N5512_io_in),
    .io_config(CBMux_IPIN22_N5512_io_config),
    .io_out(CBMux_IPIN22_N5512_io_out),
    .io_loopBreak(CBMux_IPIN22_N5512_io_loopBreak),
    .io_cnstClk(CBMux_IPIN22_N5512_io_cnstClk),
    .io_arst(CBMux_IPIN22_N5512_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN23_N5513 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN23_N5513_io_in),
    .io_config(CBMux_IPIN23_N5513_io_config),
    .io_out(CBMux_IPIN23_N5513_io_out),
    .io_loopBreak(CBMux_IPIN23_N5513_io_loopBreak),
    .io_cnstClk(CBMux_IPIN23_N5513_io_cnstClk),
    .io_arst(CBMux_IPIN23_N5513_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN24_N5514 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN24_N5514_io_in),
    .io_config(CBMux_IPIN24_N5514_io_config),
    .io_out(CBMux_IPIN24_N5514_io_out),
    .io_loopBreak(CBMux_IPIN24_N5514_io_loopBreak),
    .io_cnstClk(CBMux_IPIN24_N5514_io_cnstClk),
    .io_arst(CBMux_IPIN24_N5514_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN25_N5515 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN25_N5515_io_in),
    .io_config(CBMux_IPIN25_N5515_io_config),
    .io_out(CBMux_IPIN25_N5515_io_out),
    .io_loopBreak(CBMux_IPIN25_N5515_io_loopBreak),
    .io_cnstClk(CBMux_IPIN25_N5515_io_cnstClk),
    .io_arst(CBMux_IPIN25_N5515_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN26_N5516 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN26_N5516_io_in),
    .io_config(CBMux_IPIN26_N5516_io_config),
    .io_out(CBMux_IPIN26_N5516_io_out),
    .io_loopBreak(CBMux_IPIN26_N5516_io_loopBreak),
    .io_cnstClk(CBMux_IPIN26_N5516_io_cnstClk),
    .io_arst(CBMux_IPIN26_N5516_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN27_N5517 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN27_N5517_io_in),
    .io_config(CBMux_IPIN27_N5517_io_config),
    .io_out(CBMux_IPIN27_N5517_io_out),
    .io_loopBreak(CBMux_IPIN27_N5517_io_loopBreak),
    .io_cnstClk(CBMux_IPIN27_N5517_io_cnstClk),
    .io_arst(CBMux_IPIN27_N5517_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN28_N5518 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN28_N5518_io_in),
    .io_config(CBMux_IPIN28_N5518_io_config),
    .io_out(CBMux_IPIN28_N5518_io_out),
    .io_loopBreak(CBMux_IPIN28_N5518_io_loopBreak),
    .io_cnstClk(CBMux_IPIN28_N5518_io_cnstClk),
    .io_arst(CBMux_IPIN28_N5518_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN29_N5519 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN29_N5519_io_in),
    .io_config(CBMux_IPIN29_N5519_io_config),
    .io_out(CBMux_IPIN29_N5519_io_out),
    .io_loopBreak(CBMux_IPIN29_N5519_io_loopBreak),
    .io_cnstClk(CBMux_IPIN29_N5519_io_cnstClk),
    .io_arst(CBMux_IPIN29_N5519_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN30_N5520 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN30_N5520_io_in),
    .io_config(CBMux_IPIN30_N5520_io_config),
    .io_out(CBMux_IPIN30_N5520_io_out),
    .io_loopBreak(CBMux_IPIN30_N5520_io_loopBreak),
    .io_cnstClk(CBMux_IPIN30_N5520_io_cnstClk),
    .io_arst(CBMux_IPIN30_N5520_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN31_N5521 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN31_N5521_io_in),
    .io_config(CBMux_IPIN31_N5521_io_config),
    .io_out(CBMux_IPIN31_N5521_io_out),
    .io_loopBreak(CBMux_IPIN31_N5521_io_loopBreak),
    .io_cnstClk(CBMux_IPIN31_N5521_io_cnstClk),
    .io_arst(CBMux_IPIN31_N5521_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN32_N5522 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN32_N5522_io_in),
    .io_config(CBMux_IPIN32_N5522_io_config),
    .io_out(CBMux_IPIN32_N5522_io_out),
    .io_loopBreak(CBMux_IPIN32_N5522_io_loopBreak),
    .io_cnstClk(CBMux_IPIN32_N5522_io_cnstClk),
    .io_arst(CBMux_IPIN32_N5522_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN33_N5523 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN33_N5523_io_in),
    .io_config(CBMux_IPIN33_N5523_io_config),
    .io_out(CBMux_IPIN33_N5523_io_out),
    .io_loopBreak(CBMux_IPIN33_N5523_io_loopBreak),
    .io_cnstClk(CBMux_IPIN33_N5523_io_cnstClk),
    .io_arst(CBMux_IPIN33_N5523_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN34_N5524 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN34_N5524_io_in),
    .io_config(CBMux_IPIN34_N5524_io_config),
    .io_out(CBMux_IPIN34_N5524_io_out),
    .io_loopBreak(CBMux_IPIN34_N5524_io_loopBreak),
    .io_cnstClk(CBMux_IPIN34_N5524_io_cnstClk),
    .io_arst(CBMux_IPIN34_N5524_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN35_N5525 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN35_N5525_io_in),
    .io_config(CBMux_IPIN35_N5525_io_config),
    .io_out(CBMux_IPIN35_N5525_io_out),
    .io_loopBreak(CBMux_IPIN35_N5525_io_loopBreak),
    .io_cnstClk(CBMux_IPIN35_N5525_io_cnstClk),
    .io_arst(CBMux_IPIN35_N5525_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN36_N5526 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN36_N5526_io_in),
    .io_config(CBMux_IPIN36_N5526_io_config),
    .io_out(CBMux_IPIN36_N5526_io_out),
    .io_loopBreak(CBMux_IPIN36_N5526_io_loopBreak),
    .io_cnstClk(CBMux_IPIN36_N5526_io_cnstClk),
    .io_arst(CBMux_IPIN36_N5526_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN37_N5527 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN37_N5527_io_in),
    .io_config(CBMux_IPIN37_N5527_io_config),
    .io_out(CBMux_IPIN37_N5527_io_out),
    .io_loopBreak(CBMux_IPIN37_N5527_io_loopBreak),
    .io_cnstClk(CBMux_IPIN37_N5527_io_cnstClk),
    .io_arst(CBMux_IPIN37_N5527_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN38_N5528 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN38_N5528_io_in),
    .io_config(CBMux_IPIN38_N5528_io_config),
    .io_out(CBMux_IPIN38_N5528_io_out),
    .io_loopBreak(CBMux_IPIN38_N5528_io_loopBreak),
    .io_cnstClk(CBMux_IPIN38_N5528_io_cnstClk),
    .io_arst(CBMux_IPIN38_N5528_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN39_N5529 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN39_N5529_io_in),
    .io_config(CBMux_IPIN39_N5529_io_config),
    .io_out(CBMux_IPIN39_N5529_io_out),
    .io_loopBreak(CBMux_IPIN39_N5529_io_loopBreak),
    .io_cnstClk(CBMux_IPIN39_N5529_io_cnstClk),
    .io_arst(CBMux_IPIN39_N5529_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN40_N5530 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN40_N5530_io_in),
    .io_config(CBMux_IPIN40_N5530_io_config),
    .io_out(CBMux_IPIN40_N5530_io_out),
    .io_loopBreak(CBMux_IPIN40_N5530_io_loopBreak),
    .io_cnstClk(CBMux_IPIN40_N5530_io_cnstClk),
    .io_arst(CBMux_IPIN40_N5530_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN41_N5531 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN41_N5531_io_in),
    .io_config(CBMux_IPIN41_N5531_io_config),
    .io_out(CBMux_IPIN41_N5531_io_out),
    .io_loopBreak(CBMux_IPIN41_N5531_io_loopBreak),
    .io_cnstClk(CBMux_IPIN41_N5531_io_cnstClk),
    .io_arst(CBMux_IPIN41_N5531_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN42_N5532 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN42_N5532_io_in),
    .io_config(CBMux_IPIN42_N5532_io_config),
    .io_out(CBMux_IPIN42_N5532_io_out),
    .io_loopBreak(CBMux_IPIN42_N5532_io_loopBreak),
    .io_cnstClk(CBMux_IPIN42_N5532_io_cnstClk),
    .io_arst(CBMux_IPIN42_N5532_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN43_N5533 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN43_N5533_io_in),
    .io_config(CBMux_IPIN43_N5533_io_config),
    .io_out(CBMux_IPIN43_N5533_io_out),
    .io_loopBreak(CBMux_IPIN43_N5533_io_loopBreak),
    .io_cnstClk(CBMux_IPIN43_N5533_io_cnstClk),
    .io_arst(CBMux_IPIN43_N5533_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN44_N5534 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN44_N5534_io_in),
    .io_config(CBMux_IPIN44_N5534_io_config),
    .io_out(CBMux_IPIN44_N5534_io_out),
    .io_loopBreak(CBMux_IPIN44_N5534_io_loopBreak),
    .io_cnstClk(CBMux_IPIN44_N5534_io_cnstClk),
    .io_arst(CBMux_IPIN44_N5534_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN45_N5535 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN45_N5535_io_in),
    .io_config(CBMux_IPIN45_N5535_io_config),
    .io_out(CBMux_IPIN45_N5535_io_out),
    .io_loopBreak(CBMux_IPIN45_N5535_io_loopBreak),
    .io_cnstClk(CBMux_IPIN45_N5535_io_cnstClk),
    .io_arst(CBMux_IPIN45_N5535_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN46_N5536 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN46_N5536_io_in),
    .io_config(CBMux_IPIN46_N5536_io_config),
    .io_out(CBMux_IPIN46_N5536_io_out),
    .io_loopBreak(CBMux_IPIN46_N5536_io_loopBreak),
    .io_cnstClk(CBMux_IPIN46_N5536_io_cnstClk),
    .io_arst(CBMux_IPIN46_N5536_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN47_N5537 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN47_N5537_io_in),
    .io_config(CBMux_IPIN47_N5537_io_config),
    .io_out(CBMux_IPIN47_N5537_io_out),
    .io_loopBreak(CBMux_IPIN47_N5537_io_loopBreak),
    .io_cnstClk(CBMux_IPIN47_N5537_io_cnstClk),
    .io_arst(CBMux_IPIN47_N5537_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN48_N5538 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN48_N5538_io_in),
    .io_config(CBMux_IPIN48_N5538_io_config),
    .io_out(CBMux_IPIN48_N5538_io_out),
    .io_loopBreak(CBMux_IPIN48_N5538_io_loopBreak),
    .io_cnstClk(CBMux_IPIN48_N5538_io_cnstClk),
    .io_arst(CBMux_IPIN48_N5538_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN49_N5539 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN49_N5539_io_in),
    .io_config(CBMux_IPIN49_N5539_io_config),
    .io_out(CBMux_IPIN49_N5539_io_out),
    .io_loopBreak(CBMux_IPIN49_N5539_io_loopBreak),
    .io_cnstClk(CBMux_IPIN49_N5539_io_cnstClk),
    .io_arst(CBMux_IPIN49_N5539_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN50_N5540 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN50_N5540_io_in),
    .io_config(CBMux_IPIN50_N5540_io_config),
    .io_out(CBMux_IPIN50_N5540_io_out),
    .io_loopBreak(CBMux_IPIN50_N5540_io_loopBreak),
    .io_cnstClk(CBMux_IPIN50_N5540_io_cnstClk),
    .io_arst(CBMux_IPIN50_N5540_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN51_N5541 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN51_N5541_io_in),
    .io_config(CBMux_IPIN51_N5541_io_config),
    .io_out(CBMux_IPIN51_N5541_io_out),
    .io_loopBreak(CBMux_IPIN51_N5541_io_loopBreak),
    .io_cnstClk(CBMux_IPIN51_N5541_io_cnstClk),
    .io_arst(CBMux_IPIN51_N5541_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN52_N5542 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN52_N5542_io_in),
    .io_config(CBMux_IPIN52_N5542_io_config),
    .io_out(CBMux_IPIN52_N5542_io_out),
    .io_loopBreak(CBMux_IPIN52_N5542_io_loopBreak),
    .io_cnstClk(CBMux_IPIN52_N5542_io_cnstClk),
    .io_arst(CBMux_IPIN52_N5542_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN53_N5543 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN53_N5543_io_in),
    .io_config(CBMux_IPIN53_N5543_io_config),
    .io_out(CBMux_IPIN53_N5543_io_out),
    .io_loopBreak(CBMux_IPIN53_N5543_io_loopBreak),
    .io_cnstClk(CBMux_IPIN53_N5543_io_cnstClk),
    .io_arst(CBMux_IPIN53_N5543_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN54_N5544 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN54_N5544_io_in),
    .io_config(CBMux_IPIN54_N5544_io_config),
    .io_out(CBMux_IPIN54_N5544_io_out),
    .io_loopBreak(CBMux_IPIN54_N5544_io_loopBreak),
    .io_cnstClk(CBMux_IPIN54_N5544_io_cnstClk),
    .io_arst(CBMux_IPIN54_N5544_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN55_N5545 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN55_N5545_io_in),
    .io_config(CBMux_IPIN55_N5545_io_config),
    .io_out(CBMux_IPIN55_N5545_io_out),
    .io_loopBreak(CBMux_IPIN55_N5545_io_loopBreak),
    .io_cnstClk(CBMux_IPIN55_N5545_io_cnstClk),
    .io_arst(CBMux_IPIN55_N5545_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN56_N5546 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN56_N5546_io_in),
    .io_config(CBMux_IPIN56_N5546_io_config),
    .io_out(CBMux_IPIN56_N5546_io_out),
    .io_loopBreak(CBMux_IPIN56_N5546_io_loopBreak),
    .io_cnstClk(CBMux_IPIN56_N5546_io_cnstClk),
    .io_arst(CBMux_IPIN56_N5546_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN57_N5547 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN57_N5547_io_in),
    .io_config(CBMux_IPIN57_N5547_io_config),
    .io_out(CBMux_IPIN57_N5547_io_out),
    .io_loopBreak(CBMux_IPIN57_N5547_io_loopBreak),
    .io_cnstClk(CBMux_IPIN57_N5547_io_cnstClk),
    .io_arst(CBMux_IPIN57_N5547_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN58_N5548 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN58_N5548_io_in),
    .io_config(CBMux_IPIN58_N5548_io_config),
    .io_out(CBMux_IPIN58_N5548_io_out),
    .io_loopBreak(CBMux_IPIN58_N5548_io_loopBreak),
    .io_cnstClk(CBMux_IPIN58_N5548_io_cnstClk),
    .io_arst(CBMux_IPIN58_N5548_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN59_N5549 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN59_N5549_io_in),
    .io_config(CBMux_IPIN59_N5549_io_config),
    .io_out(CBMux_IPIN59_N5549_io_out),
    .io_loopBreak(CBMux_IPIN59_N5549_io_loopBreak),
    .io_cnstClk(CBMux_IPIN59_N5549_io_cnstClk),
    .io_arst(CBMux_IPIN59_N5549_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN60_N5550 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN60_N5550_io_in),
    .io_config(CBMux_IPIN60_N5550_io_config),
    .io_out(CBMux_IPIN60_N5550_io_out),
    .io_loopBreak(CBMux_IPIN60_N5550_io_loopBreak),
    .io_cnstClk(CBMux_IPIN60_N5550_io_cnstClk),
    .io_arst(CBMux_IPIN60_N5550_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN61_N5551 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN61_N5551_io_in),
    .io_config(CBMux_IPIN61_N5551_io_config),
    .io_out(CBMux_IPIN61_N5551_io_out),
    .io_loopBreak(CBMux_IPIN61_N5551_io_loopBreak),
    .io_cnstClk(CBMux_IPIN61_N5551_io_cnstClk),
    .io_arst(CBMux_IPIN61_N5551_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN62_N5552 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN62_N5552_io_in),
    .io_config(CBMux_IPIN62_N5552_io_config),
    .io_out(CBMux_IPIN62_N5552_io_out),
    .io_loopBreak(CBMux_IPIN62_N5552_io_loopBreak),
    .io_cnstClk(CBMux_IPIN62_N5552_io_cnstClk),
    .io_arst(CBMux_IPIN62_N5552_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN63_N5553 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN63_N5553_io_in),
    .io_config(CBMux_IPIN63_N5553_io_config),
    .io_out(CBMux_IPIN63_N5553_io_out),
    .io_loopBreak(CBMux_IPIN63_N5553_io_loopBreak),
    .io_cnstClk(CBMux_IPIN63_N5553_io_cnstClk),
    .io_arst(CBMux_IPIN63_N5553_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN64_N5554 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN64_N5554_io_in),
    .io_config(CBMux_IPIN64_N5554_io_config),
    .io_out(CBMux_IPIN64_N5554_io_out),
    .io_loopBreak(CBMux_IPIN64_N5554_io_loopBreak),
    .io_cnstClk(CBMux_IPIN64_N5554_io_cnstClk),
    .io_arst(CBMux_IPIN64_N5554_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN65_N5555 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN65_N5555_io_in),
    .io_config(CBMux_IPIN65_N5555_io_config),
    .io_out(CBMux_IPIN65_N5555_io_out),
    .io_loopBreak(CBMux_IPIN65_N5555_io_loopBreak),
    .io_cnstClk(CBMux_IPIN65_N5555_io_cnstClk),
    .io_arst(CBMux_IPIN65_N5555_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN66_N5556 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN66_N5556_io_in),
    .io_config(CBMux_IPIN66_N5556_io_config),
    .io_out(CBMux_IPIN66_N5556_io_out),
    .io_loopBreak(CBMux_IPIN66_N5556_io_loopBreak),
    .io_cnstClk(CBMux_IPIN66_N5556_io_cnstClk),
    .io_arst(CBMux_IPIN66_N5556_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN67_N5557 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN67_N5557_io_in),
    .io_config(CBMux_IPIN67_N5557_io_config),
    .io_out(CBMux_IPIN67_N5557_io_out),
    .io_loopBreak(CBMux_IPIN67_N5557_io_loopBreak),
    .io_cnstClk(CBMux_IPIN67_N5557_io_cnstClk),
    .io_arst(CBMux_IPIN67_N5557_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN68_N5558 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN68_N5558_io_in),
    .io_config(CBMux_IPIN68_N5558_io_config),
    .io_out(CBMux_IPIN68_N5558_io_out),
    .io_loopBreak(CBMux_IPIN68_N5558_io_loopBreak),
    .io_cnstClk(CBMux_IPIN68_N5558_io_cnstClk),
    .io_arst(CBMux_IPIN68_N5558_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN69_N5559 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN69_N5559_io_in),
    .io_config(CBMux_IPIN69_N5559_io_config),
    .io_out(CBMux_IPIN69_N5559_io_out),
    .io_loopBreak(CBMux_IPIN69_N5559_io_loopBreak),
    .io_cnstClk(CBMux_IPIN69_N5559_io_cnstClk),
    .io_arst(CBMux_IPIN69_N5559_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN70_N5560 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN70_N5560_io_in),
    .io_config(CBMux_IPIN70_N5560_io_config),
    .io_out(CBMux_IPIN70_N5560_io_out),
    .io_loopBreak(CBMux_IPIN70_N5560_io_loopBreak),
    .io_cnstClk(CBMux_IPIN70_N5560_io_cnstClk),
    .io_arst(CBMux_IPIN70_N5560_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN71_N5561 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN71_N5561_io_in),
    .io_config(CBMux_IPIN71_N5561_io_config),
    .io_out(CBMux_IPIN71_N5561_io_out),
    .io_loopBreak(CBMux_IPIN71_N5561_io_loopBreak),
    .io_cnstClk(CBMux_IPIN71_N5561_io_cnstClk),
    .io_arst(CBMux_IPIN71_N5561_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C5_N23993_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C5_N23993_O_3_C_6_io_in),
    .io_config(SBMux_C5_N23993_O_3_C_6_io_config),
    .io_out(SBMux_C5_N23993_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C5_N23993_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C5_N23993_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C5_N23993_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C5_N23993_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C13_N24001_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C13_N24001_O_3_C_6_io_in),
    .io_config(SBMux_C13_N24001_O_3_C_6_io_config),
    .io_out(SBMux_C13_N24001_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C13_N24001_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C13_N24001_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C13_N24001_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C13_N24001_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C21_N24009_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C21_N24009_O_3_C_6_io_in),
    .io_config(SBMux_C21_N24009_O_3_C_6_io_config),
    .io_out(SBMux_C21_N24009_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C21_N24009_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C21_N24009_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C21_N24009_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C21_N24009_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C29_N24017_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C29_N24017_O_3_C_6_io_in),
    .io_config(SBMux_C29_N24017_O_3_C_6_io_config),
    .io_out(SBMux_C29_N24017_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C29_N24017_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C29_N24017_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C29_N24017_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C29_N24017_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C37_N24025_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C37_N24025_O_3_C_6_io_in),
    .io_config(SBMux_C37_N24025_O_3_C_6_io_config),
    .io_out(SBMux_C37_N24025_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C37_N24025_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C37_N24025_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C37_N24025_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C37_N24025_O_3_C_6_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C45_N24033_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C45_N24033_O_4_C_5_io_in),
    .io_config(SBMux_C45_N24033_O_4_C_5_io_config),
    .io_out(SBMux_C45_N24033_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C45_N24033_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C45_N24033_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C45_N24033_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C45_N24033_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C53_N24041_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C53_N24041_O_4_C_5_io_in),
    .io_config(SBMux_C53_N24041_O_4_C_5_io_config),
    .io_out(SBMux_C53_N24041_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C53_N24041_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C53_N24041_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C53_N24041_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C53_N24041_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C6_SCAOptSB SBMux_C61_N24049_O_4_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C61_N24049_O_4_C_6_io_in),
    .io_config(SBMux_C61_N24049_O_4_C_6_io_config),
    .io_out(SBMux_C61_N24049_O_4_C_6_io_out),
    .io_loopBreak(SBMux_C61_N24049_O_4_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C61_N24049_O_4_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C61_N24049_O_4_C_6_io_cnstClk),
    .io_arst(SBMux_C61_N24049_O_4_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C69_N24057_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C69_N24057_O_3_C_6_io_in),
    .io_config(SBMux_C69_N24057_O_3_C_6_io_config),
    .io_out(SBMux_C69_N24057_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C69_N24057_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C69_N24057_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C69_N24057_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C69_N24057_O_3_C_6_io_arst)
  );
  MuxNInput_O0_C6_SCAOptSB SBMux_C77_N24089_O_0_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C77_N24089_O_0_C_6_io_in),
    .io_config(SBMux_C77_N24089_O_0_C_6_io_config),
    .io_out(SBMux_C77_N24089_O_0_C_6_io_out),
    .io_loopBreak(SBMux_C77_N24089_O_0_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C77_N24089_O_0_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C77_N24089_O_0_C_6_io_cnstClk),
    .io_arst(SBMux_C77_N24089_O_0_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C4_N24112_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C4_N24112_O_3_C_5_io_in),
    .io_config(SBMux_C4_N24112_O_3_C_5_io_config),
    .io_out(SBMux_C4_N24112_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C4_N24112_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C4_N24112_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C4_N24112_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C4_N24112_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C12_N24114_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C12_N24114_O_3_C_6_io_in),
    .io_config(SBMux_C12_N24114_O_3_C_6_io_config),
    .io_out(SBMux_C12_N24114_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C12_N24114_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C12_N24114_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C12_N24114_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C12_N24114_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C20_N24116_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C20_N24116_O_3_C_6_io_in),
    .io_config(SBMux_C20_N24116_O_3_C_6_io_config),
    .io_out(SBMux_C20_N24116_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C20_N24116_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C20_N24116_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C20_N24116_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C20_N24116_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C28_N24118_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C28_N24118_O_3_C_6_io_in),
    .io_config(SBMux_C28_N24118_O_3_C_6_io_config),
    .io_out(SBMux_C28_N24118_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C28_N24118_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C28_N24118_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C28_N24118_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C28_N24118_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C36_N24120_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C36_N24120_O_3_C_6_io_in),
    .io_config(SBMux_C36_N24120_O_3_C_6_io_config),
    .io_out(SBMux_C36_N24120_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C36_N24120_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C36_N24120_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C36_N24120_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C36_N24120_O_3_C_6_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C44_N24122_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C44_N24122_O_4_C_5_io_in),
    .io_config(SBMux_C44_N24122_O_4_C_5_io_config),
    .io_out(SBMux_C44_N24122_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C44_N24122_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C44_N24122_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C44_N24122_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C44_N24122_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C52_N24124_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C52_N24124_O_4_C_5_io_in),
    .io_config(SBMux_C52_N24124_O_4_C_5_io_config),
    .io_out(SBMux_C52_N24124_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C52_N24124_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C52_N24124_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C52_N24124_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C52_N24124_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C60_N24126_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C60_N24126_O_4_C_5_io_in),
    .io_config(SBMux_C60_N24126_O_4_C_5_io_config),
    .io_out(SBMux_C60_N24126_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C60_N24126_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C60_N24126_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C60_N24126_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C60_N24126_O_4_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C68_N24128_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C68_N24128_O_3_C_5_io_in),
    .io_config(SBMux_C68_N24128_O_3_C_5_io_config),
    .io_out(SBMux_C68_N24128_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C68_N24128_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C68_N24128_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C68_N24128_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C68_N24128_O_3_C_5_io_arst)
  );
  MuxNInput_O0_C4_SCAOptSB SBMux_C76_N24130_O_0_C_4 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C76_N24130_O_0_C_4_io_in),
    .io_config(SBMux_C76_N24130_O_0_C_4_io_config),
    .io_out(SBMux_C76_N24130_O_0_C_4_io_out),
    .io_loopBreak(SBMux_C76_N24130_O_0_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C76_N24130_O_0_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C76_N24130_O_0_C_4_io_cnstClk),
    .io_arst(SBMux_C76_N24130_O_0_C_4_io_arst)
  );
  MuxNInput_O4_C6_SCAOptSB SBMux_C5_N27119_O_4_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C5_N27119_O_4_C_6_io_in),
    .io_config(SBMux_C5_N27119_O_4_C_6_io_config),
    .io_out(SBMux_C5_N27119_O_4_C_6_io_out),
    .io_loopBreak(SBMux_C5_N27119_O_4_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C5_N27119_O_4_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C5_N27119_O_4_C_6_io_cnstClk),
    .io_arst(SBMux_C5_N27119_O_4_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C13_N27127_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C13_N27127_O_3_C_6_io_in),
    .io_config(SBMux_C13_N27127_O_3_C_6_io_config),
    .io_out(SBMux_C13_N27127_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C13_N27127_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C13_N27127_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C13_N27127_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C13_N27127_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C21_N27135_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C21_N27135_O_3_C_6_io_in),
    .io_config(SBMux_C21_N27135_O_3_C_6_io_config),
    .io_out(SBMux_C21_N27135_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C21_N27135_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C21_N27135_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C21_N27135_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C21_N27135_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C29_N27143_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C29_N27143_O_3_C_5_io_in),
    .io_config(SBMux_C29_N27143_O_3_C_5_io_config),
    .io_out(SBMux_C29_N27143_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C29_N27143_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C29_N27143_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C29_N27143_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C29_N27143_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C37_N27151_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C37_N27151_O_3_C_5_io_in),
    .io_config(SBMux_C37_N27151_O_3_C_5_io_config),
    .io_out(SBMux_C37_N27151_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C37_N27151_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C37_N27151_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C37_N27151_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C37_N27151_O_3_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C45_N27159_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C45_N27159_O_4_C_5_io_in),
    .io_config(SBMux_C45_N27159_O_4_C_5_io_config),
    .io_out(SBMux_C45_N27159_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C45_N27159_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C45_N27159_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C45_N27159_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C45_N27159_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C53_N27167_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C53_N27167_O_4_C_5_io_in),
    .io_config(SBMux_C53_N27167_O_4_C_5_io_config),
    .io_out(SBMux_C53_N27167_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C53_N27167_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C53_N27167_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C53_N27167_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C53_N27167_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C61_N27175_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C61_N27175_O_4_C_5_io_in),
    .io_config(SBMux_C61_N27175_O_4_C_5_io_config),
    .io_out(SBMux_C61_N27175_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C61_N27175_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C61_N27175_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C61_N27175_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C61_N27175_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C69_N27183_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C69_N27183_O_4_C_5_io_in),
    .io_config(SBMux_C69_N27183_O_4_C_5_io_config),
    .io_out(SBMux_C69_N27183_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C69_N27183_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C69_N27183_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C69_N27183_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C69_N27183_O_4_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C77_N27215_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C77_N27215_O_3_C_5_io_in),
    .io_config(SBMux_C77_N27215_O_3_C_5_io_config),
    .io_out(SBMux_C77_N27215_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C77_N27215_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C77_N27215_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C77_N27215_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C77_N27215_O_3_C_5_io_arst)
  );
  MuxNInput_O4_C7_SCAOptSB SBMux_C4_N27238_O_4_C_7 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C4_N27238_O_4_C_7_io_in),
    .io_config(SBMux_C4_N27238_O_4_C_7_io_config),
    .io_out(SBMux_C4_N27238_O_4_C_7_io_out),
    .io_loopBreak(SBMux_C4_N27238_O_4_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C4_N27238_O_4_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C4_N27238_O_4_C_7_io_cnstClk),
    .io_arst(SBMux_C4_N27238_O_4_C_7_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C12_N27240_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C12_N27240_O_3_C_6_io_in),
    .io_config(SBMux_C12_N27240_O_3_C_6_io_config),
    .io_out(SBMux_C12_N27240_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C12_N27240_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C12_N27240_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C12_N27240_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C12_N27240_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C20_N27242_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C20_N27242_O_3_C_6_io_in),
    .io_config(SBMux_C20_N27242_O_3_C_6_io_config),
    .io_out(SBMux_C20_N27242_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C20_N27242_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C20_N27242_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C20_N27242_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C20_N27242_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C28_N27244_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C28_N27244_O_3_C_5_io_in),
    .io_config(SBMux_C28_N27244_O_3_C_5_io_config),
    .io_out(SBMux_C28_N27244_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C28_N27244_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C28_N27244_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C28_N27244_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C28_N27244_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C36_N27246_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C36_N27246_O_3_C_5_io_in),
    .io_config(SBMux_C36_N27246_O_3_C_5_io_config),
    .io_out(SBMux_C36_N27246_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C36_N27246_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C36_N27246_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C36_N27246_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C36_N27246_O_3_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C44_N27248_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C44_N27248_O_4_C_5_io_in),
    .io_config(SBMux_C44_N27248_O_4_C_5_io_config),
    .io_out(SBMux_C44_N27248_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C44_N27248_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C44_N27248_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C44_N27248_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C44_N27248_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C52_N27250_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C52_N27250_O_4_C_5_io_in),
    .io_config(SBMux_C52_N27250_O_4_C_5_io_config),
    .io_out(SBMux_C52_N27250_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C52_N27250_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C52_N27250_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C52_N27250_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C52_N27250_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C6_SCAOptSB SBMux_C60_N27252_O_4_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C60_N27252_O_4_C_6_io_in),
    .io_config(SBMux_C60_N27252_O_4_C_6_io_config),
    .io_out(SBMux_C60_N27252_O_4_C_6_io_out),
    .io_loopBreak(SBMux_C60_N27252_O_4_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C60_N27252_O_4_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C60_N27252_O_4_C_6_io_cnstClk),
    .io_arst(SBMux_C60_N27252_O_4_C_6_io_arst)
  );
  MuxNInput_O4_C6_SCAOptSB SBMux_C68_N27254_O_4_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C68_N27254_O_4_C_6_io_in),
    .io_config(SBMux_C68_N27254_O_4_C_6_io_config),
    .io_out(SBMux_C68_N27254_O_4_C_6_io_out),
    .io_loopBreak(SBMux_C68_N27254_O_4_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C68_N27254_O_4_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C68_N27254_O_4_C_6_io_cnstClk),
    .io_arst(SBMux_C68_N27254_O_4_C_6_io_arst)
  );
  MuxNInput_O3_C7_SCAOptSB SBMux_C76_N27256_O_3_C_7 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C76_N27256_O_3_C_7_io_in),
    .io_config(SBMux_C76_N27256_O_3_C_7_io_config),
    .io_out(SBMux_C76_N27256_O_3_C_7_io_out),
    .io_loopBreak(SBMux_C76_N27256_O_3_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C76_N27256_O_3_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C76_N27256_O_3_C_7_io_cnstClk),
    .io_arst(SBMux_C76_N27256_O_3_C_7_io_arst)
  );
  assign OUT_OPIN_N5581_91 = logicBlock_OPIN_91; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5603_113 = logicBlock_OPIN_113; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5572_82 = logicBlock_OPIN_82; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5610_120 = logicBlock_OPIN_120; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N27159_45 = SBMux_C45_N27159_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24009_21 = SBMux_C21_N24009_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5577_87 = logicBlock_OPIN_87; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N27240_12 = SBMux_C12_N27240_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N27151_37 = SBMux_C37_N27151_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5600_110 = logicBlock_OPIN_110; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5566_76 = logicBlock_OPIN_76; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N27254_68 = SBMux_C68_N27254_O_4_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N27143_29 = SBMux_C29_N27143_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5595_105 = logicBlock_OPIN_105; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24120_36 = SBMux_C36_N24120_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N27244_28 = SBMux_C28_N27244_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5601_111 = logicBlock_OPIN_111; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N27242_20 = SBMux_C20_N27242_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N27119_5 = SBMux_C5_N27119_O_4_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5609_119 = logicBlock_OPIN_119; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5588_98 = logicBlock_OPIN_98; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24126_60 = SBMux_C60_N24126_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5604_114 = logicBlock_OPIN_114; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24033_45 = SBMux_C45_N24033_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N27175_61 = SBMux_C61_N27175_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N27250_52 = SBMux_C52_N27250_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24112_4 = SBMux_C4_N24112_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24057_69 = SBMux_C69_N24057_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24130_76 = SBMux_C76_N24130_O_0_C_4_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N27252_60 = SBMux_C60_N27252_O_4_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5585_95 = logicBlock_OPIN_95; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N27246_36 = SBMux_C36_N27246_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5586_96 = logicBlock_OPIN_96; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24041_53 = SBMux_C53_N24041_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5568_78 = logicBlock_OPIN_78; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5592_102 = logicBlock_OPIN_102; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5583_93 = logicBlock_OPIN_93; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5605_115 = logicBlock_OPIN_115; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5608_118 = logicBlock_OPIN_118; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24118_28 = SBMux_C28_N24118_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5596_106 = logicBlock_OPIN_106; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5571_81 = logicBlock_OPIN_81; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5563_73 = logicBlock_OPIN_73; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5576_86 = logicBlock_OPIN_86; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5582_92 = logicBlock_OPIN_92; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24128_68 = SBMux_C68_N24128_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5573_83 = logicBlock_OPIN_83; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24017_29 = SBMux_C29_N24017_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5580_90 = logicBlock_OPIN_90; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5606_116 = logicBlock_OPIN_116; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24124_52 = SBMux_C52_N24124_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5598_108 = logicBlock_OPIN_108; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24049_61 = SBMux_C61_N24049_O_4_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5589_99 = logicBlock_OPIN_99; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5567_77 = logicBlock_OPIN_77; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5591_101 = logicBlock_OPIN_101; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5597_107 = logicBlock_OPIN_107; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5569_79 = logicBlock_OPIN_79; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N27238_4 = SBMux_C4_N27238_O_4_C_7_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5570_80 = logicBlock_OPIN_80; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N27183_69 = SBMux_C69_N27183_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5593_103 = logicBlock_OPIN_103; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5574_84 = logicBlock_OPIN_84; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24114_12 = SBMux_C12_N24114_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5575_85 = logicBlock_OPIN_85; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5599_109 = logicBlock_OPIN_109; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5584_94 = logicBlock_OPIN_94; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5578_88 = logicBlock_OPIN_88; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5579_89 = logicBlock_OPIN_89; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24025_37 = SBMux_C37_N24025_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5565_75 = logicBlock_OPIN_75; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5564_74 = logicBlock_OPIN_74; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N5587_97 = logicBlock_OPIN_97; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N27215_77 = SBMux_C77_N27215_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5607_117 = logicBlock_OPIN_117; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N27256_76 = SBMux_C76_N27256_O_3_C_7_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N23993_5 = SBMux_C5_N23993_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5594_104 = logicBlock_OPIN_104; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N27135_21 = SBMux_C21_N27135_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N27167_53 = SBMux_C53_N27167_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24001_13 = SBMux_C13_N24001_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N27127_13 = SBMux_C13_N27127_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5590_100 = logicBlock_OPIN_100; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24116_20 = SBMux_C20_N24116_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24122_44 = SBMux_C44_N24122_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N27248_44 = SBMux_C44_N27248_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N5602_112 = logicBlock_OPIN_112; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24089_77 = SBMux_C77_N24089_O_0_C_6_io_out; // @[TileFull.scala 138:23]
  assign ioConf_confOut = configBlock_ioBundle_confOut; // @[TileFull.scala 73:12]
  assign ioConf_scan_out = configBlock_ioBundle_scan_out; // @[TileFull.scala 73:12]
  assign logicBlock_IPIN_0 = CBMux_IPIN0_N5490_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_1 = CBMux_IPIN1_N5491_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_2 = CBMux_IPIN2_N5492_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_3 = CBMux_IPIN3_N5493_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_4 = CBMux_IPIN4_N5494_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_5 = CBMux_IPIN5_N5495_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_6 = CBMux_IPIN6_N5496_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_7 = CBMux_IPIN7_N5497_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_8 = CBMux_IPIN8_N5498_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_9 = CBMux_IPIN9_N5499_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_10 = CBMux_IPIN10_N5500_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_11 = CBMux_IPIN11_N5501_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_12 = CBMux_IPIN12_N5502_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_13 = CBMux_IPIN13_N5503_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_14 = CBMux_IPIN14_N5504_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_15 = CBMux_IPIN15_N5505_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_16 = CBMux_IPIN16_N5506_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_17 = CBMux_IPIN17_N5507_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_18 = CBMux_IPIN18_N5508_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_19 = CBMux_IPIN19_N5509_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_20 = CBMux_IPIN20_N5510_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_21 = CBMux_IPIN21_N5511_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_22 = CBMux_IPIN22_N5512_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_23 = CBMux_IPIN23_N5513_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_24 = CBMux_IPIN24_N5514_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_25 = CBMux_IPIN25_N5515_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_26 = CBMux_IPIN26_N5516_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_27 = CBMux_IPIN27_N5517_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_28 = CBMux_IPIN28_N5518_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_29 = CBMux_IPIN29_N5519_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_30 = CBMux_IPIN30_N5520_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_31 = CBMux_IPIN31_N5521_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_32 = CBMux_IPIN32_N5522_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_33 = CBMux_IPIN33_N5523_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_34 = CBMux_IPIN34_N5524_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_35 = CBMux_IPIN35_N5525_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_36 = CBMux_IPIN36_N5526_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_37 = CBMux_IPIN37_N5527_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_38 = CBMux_IPIN38_N5528_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_39 = CBMux_IPIN39_N5529_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_40 = CBMux_IPIN40_N5530_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_41 = CBMux_IPIN41_N5531_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_42 = CBMux_IPIN42_N5532_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_43 = CBMux_IPIN43_N5533_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_44 = CBMux_IPIN44_N5534_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_45 = CBMux_IPIN45_N5535_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_46 = CBMux_IPIN46_N5536_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_47 = CBMux_IPIN47_N5537_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_48 = CBMux_IPIN48_N5538_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_49 = CBMux_IPIN49_N5539_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_50 = CBMux_IPIN50_N5540_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_51 = CBMux_IPIN51_N5541_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_52 = CBMux_IPIN52_N5542_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_53 = CBMux_IPIN53_N5543_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_54 = CBMux_IPIN54_N5544_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_55 = CBMux_IPIN55_N5545_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_56 = CBMux_IPIN56_N5546_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_57 = CBMux_IPIN57_N5547_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_58 = CBMux_IPIN58_N5548_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_59 = CBMux_IPIN59_N5549_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_60 = CBMux_IPIN60_N5550_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_61 = CBMux_IPIN61_N5551_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_62 = CBMux_IPIN62_N5552_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_63 = CBMux_IPIN63_N5553_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_64 = CBMux_IPIN64_N5554_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_65 = CBMux_IPIN65_N5555_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_66 = CBMux_IPIN66_N5556_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_67 = CBMux_IPIN67_N5557_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_68 = CBMux_IPIN68_N5558_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_69 = CBMux_IPIN69_N5559_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_70 = CBMux_IPIN70_N5560_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_71 = CBMux_IPIN71_N5561_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_clock = clock; // @[TileFull.scala 192:26]
  assign logicBlock_reset = reset; // @[TileFull.scala 193:26]
  assign logicBlock_configBits = configBlock_ioBundle_confOut[193:0]; // @[TileFull.scala 191:31]
  assign logicBlock_gndLBouts = ctrlSignals_gndBlkOuts; // @[TileFull.scala 189:30]
  assign configBlock_clock = ctrlSignals_confClock; // @[TileFull.scala 74:27]
  assign configBlock_ioBundle_scan_in = ioConf_scan_in; // @[TileFull.scala 73:12]
  assign configBlock_ioBundle_scan_en = ioConf_scan_en; // @[TileFull.scala 73:12]
  assign CBMux_IPIN0_N5490_io_in = {CBMux_IPIN0_N5490_io_in_hi,CBMux_IPIN0_N5490_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN0_N5490_io_config = configBlock_ioBundle_confOut[163:160]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN0_N5490_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN0_N5490_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN0_N5490_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN1_N5491_io_in = {CBMux_IPIN1_N5491_io_in_hi,CBMux_IPIN1_N5491_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN1_N5491_io_config = configBlock_ioBundle_confOut[167:164]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN1_N5491_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN1_N5491_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN1_N5491_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN2_N5492_io_in = {CBMux_IPIN2_N5492_io_in_hi,CBMux_IPIN2_N5492_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN2_N5492_io_config = configBlock_ioBundle_confOut[171:168]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN2_N5492_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN2_N5492_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN2_N5492_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN3_N5493_io_in = {CBMux_IPIN3_N5493_io_in_hi,CBMux_IPIN3_N5493_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN3_N5493_io_config = configBlock_ioBundle_confOut[176:172]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN3_N5493_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN3_N5493_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN3_N5493_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN4_N5494_io_in = {CBMux_IPIN4_N5494_io_in_hi,CBMux_IPIN4_N5494_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN4_N5494_io_config = configBlock_ioBundle_confOut[180:177]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN4_N5494_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN4_N5494_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN4_N5494_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN5_N5495_io_in = {CBMux_IPIN5_N5495_io_in_hi,CBMux_IPIN5_N5495_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN5_N5495_io_config = configBlock_ioBundle_confOut[184:181]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN5_N5495_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN5_N5495_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN5_N5495_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN6_N5496_io_in = {CBMux_IPIN6_N5496_io_in_hi,CBMux_IPIN6_N5496_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN6_N5496_io_config = configBlock_ioBundle_confOut[188:185]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN6_N5496_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN6_N5496_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN6_N5496_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN7_N5497_io_in = {CBMux_IPIN7_N5497_io_in_hi,CBMux_IPIN7_N5497_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN7_N5497_io_config = configBlock_ioBundle_confOut[192:189]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN7_N5497_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN7_N5497_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN7_N5497_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN8_N5498_io_in = {CBMux_IPIN8_N5498_io_in_hi,CBMux_IPIN8_N5498_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN8_N5498_io_config = configBlock_ioBundle_confOut[196:193]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN8_N5498_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN8_N5498_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN8_N5498_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN9_N5499_io_in = {CBMux_IPIN9_N5499_io_in_hi,CBMux_IPIN9_N5499_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN9_N5499_io_config = configBlock_ioBundle_confOut[200:197]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN9_N5499_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN9_N5499_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN9_N5499_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN10_N5500_io_in = {CBMux_IPIN10_N5500_io_in_hi,CBMux_IPIN10_N5500_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN10_N5500_io_config = configBlock_ioBundle_confOut[204:201]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN10_N5500_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN10_N5500_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN10_N5500_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN11_N5501_io_in = {CBMux_IPIN11_N5501_io_in_hi,CBMux_IPIN11_N5501_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN11_N5501_io_config = configBlock_ioBundle_confOut[208:205]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN11_N5501_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN11_N5501_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN11_N5501_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN12_N5502_io_in = {CBMux_IPIN12_N5502_io_in_hi,CBMux_IPIN12_N5502_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN12_N5502_io_config = configBlock_ioBundle_confOut[212:209]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN12_N5502_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN12_N5502_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN12_N5502_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN13_N5503_io_in = {CBMux_IPIN13_N5503_io_in_hi,CBMux_IPIN13_N5503_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN13_N5503_io_config = configBlock_ioBundle_confOut[216:213]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN13_N5503_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN13_N5503_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN13_N5503_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN14_N5504_io_in = {CBMux_IPIN2_N5492_io_in_hi,CBMux_IPIN14_N5504_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN14_N5504_io_config = configBlock_ioBundle_confOut[220:217]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN14_N5504_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN14_N5504_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN14_N5504_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN15_N5505_io_in = {CBMux_IPIN15_N5505_io_in_hi,CBMux_IPIN15_N5505_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN15_N5505_io_config = configBlock_ioBundle_confOut[224:221]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN15_N5505_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN15_N5505_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN15_N5505_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN16_N5506_io_in = {CBMux_IPIN16_N5506_io_in_hi,CBMux_IPIN16_N5506_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN16_N5506_io_config = configBlock_ioBundle_confOut[228:225]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN16_N5506_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN16_N5506_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN16_N5506_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN17_N5507_io_in = {CBMux_IPIN17_N5507_io_in_hi,CBMux_IPIN17_N5507_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN17_N5507_io_config = configBlock_ioBundle_confOut[232:229]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN17_N5507_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN17_N5507_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN17_N5507_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN18_N5508_io_in = {CBMux_IPIN18_N5508_io_in_hi,CBMux_IPIN18_N5508_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN18_N5508_io_config = configBlock_ioBundle_confOut[236:233]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN18_N5508_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN18_N5508_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN18_N5508_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN19_N5509_io_in = {CBMux_IPIN19_N5509_io_in_hi,CBMux_IPIN19_N5509_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN19_N5509_io_config = configBlock_ioBundle_confOut[240:237]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN19_N5509_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN19_N5509_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN19_N5509_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN20_N5510_io_in = {CBMux_IPIN20_N5510_io_in_hi,CBMux_IPIN20_N5510_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN20_N5510_io_config = configBlock_ioBundle_confOut[244:241]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN20_N5510_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN20_N5510_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN20_N5510_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN21_N5511_io_in = {CBMux_IPIN21_N5511_io_in_hi,CBMux_IPIN21_N5511_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN21_N5511_io_config = configBlock_ioBundle_confOut[248:245]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN21_N5511_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN21_N5511_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN21_N5511_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN22_N5512_io_in = {CBMux_IPIN16_N5506_io_in_hi,CBMux_IPIN22_N5512_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN22_N5512_io_config = configBlock_ioBundle_confOut[252:249]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN22_N5512_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN22_N5512_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN22_N5512_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN23_N5513_io_in = {CBMux_IPIN23_N5513_io_in_hi,CBMux_IPIN23_N5513_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN23_N5513_io_config = configBlock_ioBundle_confOut[256:253]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN23_N5513_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN23_N5513_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN23_N5513_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN24_N5514_io_in = {CBMux_IPIN24_N5514_io_in_hi,CBMux_IPIN24_N5514_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN24_N5514_io_config = configBlock_ioBundle_confOut[260:257]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN24_N5514_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN24_N5514_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN24_N5514_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN25_N5515_io_in = {CBMux_IPIN25_N5515_io_in_hi,CBMux_IPIN25_N5515_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN25_N5515_io_config = configBlock_ioBundle_confOut[264:261]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN25_N5515_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN25_N5515_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN25_N5515_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN26_N5516_io_in = {CBMux_IPIN26_N5516_io_in_hi,CBMux_IPIN26_N5516_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN26_N5516_io_config = configBlock_ioBundle_confOut[268:265]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN26_N5516_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN26_N5516_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN26_N5516_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN27_N5517_io_in = {CBMux_IPIN21_N5511_io_in_hi,CBMux_IPIN27_N5517_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN27_N5517_io_config = configBlock_ioBundle_confOut[272:269]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN27_N5517_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN27_N5517_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN27_N5517_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN28_N5518_io_in = {CBMux_IPIN28_N5518_io_in_hi,CBMux_IPIN22_N5512_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN28_N5518_io_config = configBlock_ioBundle_confOut[276:273]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN28_N5518_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN28_N5518_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN28_N5518_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN29_N5519_io_in = {CBMux_IPIN29_N5519_io_in_hi,CBMux_IPIN29_N5519_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN29_N5519_io_config = configBlock_ioBundle_confOut[280:277]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN29_N5519_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN29_N5519_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN29_N5519_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN30_N5520_io_in = {CBMux_IPIN18_N5508_io_in_hi,CBMux_IPIN30_N5520_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN30_N5520_io_config = configBlock_ioBundle_confOut[284:281]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN30_N5520_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN30_N5520_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN30_N5520_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN31_N5521_io_in = {CBMux_IPIN31_N5521_io_in_hi,CBMux_IPIN31_N5521_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN31_N5521_io_config = configBlock_ioBundle_confOut[288:285]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN31_N5521_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN31_N5521_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN31_N5521_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN32_N5522_io_in = {CBMux_IPIN32_N5522_io_in_hi,CBMux_IPIN32_N5522_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN32_N5522_io_config = configBlock_ioBundle_confOut[292:289]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN32_N5522_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN32_N5522_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN32_N5522_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN33_N5523_io_in = {CBMux_IPIN33_N5523_io_in_hi,CBMux_IPIN27_N5517_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN33_N5523_io_config = configBlock_ioBundle_confOut[296:293]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN33_N5523_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN33_N5523_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN33_N5523_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN34_N5524_io_in = {CBMux_IPIN34_N5524_io_in_hi,CBMux_IPIN34_N5524_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN34_N5524_io_config = configBlock_ioBundle_confOut[300:297]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN34_N5524_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN34_N5524_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN34_N5524_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN35_N5525_io_in = {CBMux_IPIN34_N5524_io_in_hi,CBMux_IPIN34_N5524_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN35_N5525_io_config = configBlock_ioBundle_confOut[304:301]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN35_N5525_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN35_N5525_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN35_N5525_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN36_N5526_io_in = {CBMux_IPIN36_N5526_io_in_hi,CBMux_IPIN36_N5526_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN36_N5526_io_config = configBlock_ioBundle_confOut[308:305]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN36_N5526_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN36_N5526_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN36_N5526_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN37_N5527_io_in = {CBMux_IPIN37_N5527_io_in_hi,CBMux_IPIN37_N5527_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN37_N5527_io_config = configBlock_ioBundle_confOut[312:309]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN37_N5527_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN37_N5527_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN37_N5527_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN38_N5528_io_in = {CBMux_IPIN20_N5510_io_in_hi,CBMux_IPIN20_N5510_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN38_N5528_io_config = configBlock_ioBundle_confOut[316:313]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN38_N5528_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN38_N5528_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN38_N5528_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN39_N5529_io_in = {CBMux_IPIN33_N5523_io_in_hi,CBMux_IPIN27_N5517_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN39_N5529_io_config = configBlock_ioBundle_confOut[320:317]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN39_N5529_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN39_N5529_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN39_N5529_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN40_N5530_io_in = IN_OPIN_N5823_89; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN40_N5530_io_config = configBlock_ioBundle_confOut[321]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN40_N5530_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN40_N5530_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN40_N5530_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN41_N5531_io_in = IN_OPIN_N5824_90; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN41_N5531_io_config = configBlock_ioBundle_confOut[322]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN41_N5531_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN41_N5531_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN41_N5531_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN42_N5532_io_in = IN_OPIN_N5825_91; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN42_N5532_io_config = configBlock_ioBundle_confOut[323]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN42_N5532_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN42_N5532_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN42_N5532_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN43_N5533_io_in = IN_OPIN_N5826_92; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN43_N5533_io_config = configBlock_ioBundle_confOut[324]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN43_N5533_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN43_N5533_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN43_N5533_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN44_N5534_io_in = IN_OPIN_N5827_93; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN44_N5534_io_config = configBlock_ioBundle_confOut[325]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN44_N5534_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN44_N5534_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN44_N5534_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN45_N5535_io_in = IN_OPIN_N5828_94; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN45_N5535_io_config = configBlock_ioBundle_confOut[326]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN45_N5535_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN45_N5535_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN45_N5535_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN46_N5536_io_in = IN_OPIN_N5829_95; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN46_N5536_io_config = configBlock_ioBundle_confOut[327]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN46_N5536_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN46_N5536_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN46_N5536_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN47_N5537_io_in = IN_OPIN_N5830_96; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN47_N5537_io_config = configBlock_ioBundle_confOut[328]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN47_N5537_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN47_N5537_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN47_N5537_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN48_N5538_io_in = IN_OPIN_N5831_97; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN48_N5538_io_config = configBlock_ioBundle_confOut[329]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN48_N5538_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN48_N5538_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN48_N5538_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN49_N5539_io_in = IN_OPIN_N5832_98; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN49_N5539_io_config = configBlock_ioBundle_confOut[330]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN49_N5539_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN49_N5539_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN49_N5539_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN50_N5540_io_in = IN_OPIN_N5833_99; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN50_N5540_io_config = configBlock_ioBundle_confOut[331]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN50_N5540_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN50_N5540_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN50_N5540_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN51_N5541_io_in = IN_OPIN_N5834_100; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN51_N5541_io_config = configBlock_ioBundle_confOut[332]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN51_N5541_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN51_N5541_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN51_N5541_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN52_N5542_io_in = IN_OPIN_N5835_101; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN52_N5542_io_config = configBlock_ioBundle_confOut[333]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN52_N5542_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN52_N5542_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN52_N5542_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN53_N5543_io_in = IN_OPIN_N5836_102; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN53_N5543_io_config = configBlock_ioBundle_confOut[334]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN53_N5543_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN53_N5543_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN53_N5543_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN54_N5544_io_in = IN_OPIN_N5837_103; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN54_N5544_io_config = configBlock_ioBundle_confOut[335]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN54_N5544_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN54_N5544_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN54_N5544_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN55_N5545_io_in = IN_OPIN_N5838_104; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN55_N5545_io_config = configBlock_ioBundle_confOut[336]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN55_N5545_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN55_N5545_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN55_N5545_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN56_N5546_io_in = IN_OPIN_N5839_105; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN56_N5546_io_config = configBlock_ioBundle_confOut[337]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN56_N5546_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN56_N5546_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN56_N5546_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN57_N5547_io_in = IN_OPIN_N5840_106; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN57_N5547_io_config = configBlock_ioBundle_confOut[338]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN57_N5547_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN57_N5547_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN57_N5547_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN58_N5548_io_in = IN_OPIN_N5841_107; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN58_N5548_io_config = configBlock_ioBundle_confOut[339]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN58_N5548_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN58_N5548_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN58_N5548_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN59_N5549_io_in = IN_OPIN_N5842_108; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN59_N5549_io_config = configBlock_ioBundle_confOut[340]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN59_N5549_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN59_N5549_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN59_N5549_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN60_N5550_io_in = IN_OPIN_N5843_109; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN60_N5550_io_config = configBlock_ioBundle_confOut[341]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN60_N5550_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN60_N5550_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN60_N5550_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN61_N5551_io_in = IN_OPIN_N5844_110; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN61_N5551_io_config = configBlock_ioBundle_confOut[342]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN61_N5551_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN61_N5551_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN61_N5551_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN62_N5552_io_in = IN_OPIN_N5845_111; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN62_N5552_io_config = configBlock_ioBundle_confOut[343]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN62_N5552_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN62_N5552_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN62_N5552_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN63_N5553_io_in = IN_OPIN_N5846_112; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN63_N5553_io_config = configBlock_ioBundle_confOut[344]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN63_N5553_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN63_N5553_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN63_N5553_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN64_N5554_io_in = IN_OPIN_N5847_113; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN64_N5554_io_config = configBlock_ioBundle_confOut[345]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN64_N5554_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN64_N5554_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN64_N5554_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN65_N5555_io_in = IN_OPIN_N5848_114; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN65_N5555_io_config = configBlock_ioBundle_confOut[346]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN65_N5555_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN65_N5555_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN65_N5555_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN66_N5556_io_in = IN_OPIN_N5849_115; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN66_N5556_io_config = configBlock_ioBundle_confOut[347]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN66_N5556_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN66_N5556_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN66_N5556_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN67_N5557_io_in = IN_OPIN_N5850_116; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN67_N5557_io_config = configBlock_ioBundle_confOut[348]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN67_N5557_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN67_N5557_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN67_N5557_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN68_N5558_io_in = IN_OPIN_N5851_117; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN68_N5558_io_config = configBlock_ioBundle_confOut[349]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN68_N5558_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN68_N5558_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN68_N5558_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN69_N5559_io_in = IN_OPIN_N5852_118; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN69_N5559_io_config = configBlock_ioBundle_confOut[350]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN69_N5559_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN69_N5559_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN69_N5559_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN70_N5560_io_in = IN_OPIN_N5853_119; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN70_N5560_io_config = configBlock_ioBundle_confOut[351]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN70_N5560_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN70_N5560_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN70_N5560_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN71_N5561_io_in = IN_OPIN_N5854_120; // @[TileFull.scala 161:{37,37}]
  assign CBMux_IPIN71_N5561_io_config = configBlock_ioBundle_confOut[352]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN71_N5561_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN71_N5561_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN71_N5561_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign SBMux_C5_N23993_O_3_C_6_io_in = {SBMux_C5_N23993_O_3_C_6_io_in_hi,SBMux_C5_N23993_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C5_N23993_O_3_C_6_io_config = configBlock_ioBundle_confOut[356:353]; // @[TileFull.scala 142:60]
  assign SBMux_C5_N23993_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C5_N23993_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C5_N23993_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C5_N23993_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C13_N24001_O_3_C_6_io_in = {SBMux_C13_N24001_O_3_C_6_io_in_hi,SBMux_C13_N24001_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C13_N24001_O_3_C_6_io_config = configBlock_ioBundle_confOut[360:357]; // @[TileFull.scala 142:60]
  assign SBMux_C13_N24001_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C13_N24001_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C13_N24001_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C13_N24001_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C21_N24009_O_3_C_6_io_in = {SBMux_C21_N24009_O_3_C_6_io_in_hi,SBMux_C21_N24009_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C21_N24009_O_3_C_6_io_config = configBlock_ioBundle_confOut[364:361]; // @[TileFull.scala 142:60]
  assign SBMux_C21_N24009_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C21_N24009_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C21_N24009_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C21_N24009_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C29_N24017_O_3_C_6_io_in = {SBMux_C29_N24017_O_3_C_6_io_in_hi,SBMux_C29_N24017_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C29_N24017_O_3_C_6_io_config = configBlock_ioBundle_confOut[368:365]; // @[TileFull.scala 142:60]
  assign SBMux_C29_N24017_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C29_N24017_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C29_N24017_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C29_N24017_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C37_N24025_O_3_C_6_io_in = {SBMux_C37_N24025_O_3_C_6_io_in_hi,SBMux_C37_N24025_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C37_N24025_O_3_C_6_io_config = configBlock_ioBundle_confOut[372:369]; // @[TileFull.scala 142:60]
  assign SBMux_C37_N24025_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C37_N24025_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C37_N24025_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C37_N24025_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C45_N24033_O_4_C_5_io_in = {SBMux_C45_N24033_O_4_C_5_io_in_hi,SBMux_C45_N24033_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C45_N24033_O_4_C_5_io_config = configBlock_ioBundle_confOut[376:373]; // @[TileFull.scala 142:60]
  assign SBMux_C45_N24033_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C45_N24033_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C45_N24033_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C45_N24033_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C53_N24041_O_4_C_5_io_in = {SBMux_C53_N24041_O_4_C_5_io_in_hi,SBMux_C45_N24033_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C53_N24041_O_4_C_5_io_config = configBlock_ioBundle_confOut[380:377]; // @[TileFull.scala 142:60]
  assign SBMux_C53_N24041_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C53_N24041_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C53_N24041_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C53_N24041_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C61_N24049_O_4_C_6_io_in = {SBMux_C61_N24049_O_4_C_6_io_in_hi,SBMux_C61_N24049_O_4_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C61_N24049_O_4_C_6_io_config = configBlock_ioBundle_confOut[384:381]; // @[TileFull.scala 142:60]
  assign SBMux_C61_N24049_O_4_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C61_N24049_O_4_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C61_N24049_O_4_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C61_N24049_O_4_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C69_N24057_O_3_C_6_io_in = {SBMux_C69_N24057_O_3_C_6_io_in_hi,SBMux_C69_N24057_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C69_N24057_O_3_C_6_io_config = configBlock_ioBundle_confOut[388:385]; // @[TileFull.scala 142:60]
  assign SBMux_C69_N24057_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C69_N24057_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C69_N24057_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C69_N24057_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C77_N24089_O_0_C_6_io_in = {SBMux_C77_N24089_O_0_C_6_io_in_hi,SBMux_C77_N24089_O_0_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C77_N24089_O_0_C_6_io_config = configBlock_ioBundle_confOut[392:389]; // @[TileFull.scala 142:60]
  assign SBMux_C77_N24089_O_0_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C77_N24089_O_0_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C77_N24089_O_0_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C77_N24089_O_0_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C4_N24112_O_3_C_5_io_in = {SBMux_C4_N24112_O_3_C_5_io_in_hi,SBMux_C4_N24112_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C4_N24112_O_3_C_5_io_config = configBlock_ioBundle_confOut[396:393]; // @[TileFull.scala 142:60]
  assign SBMux_C4_N24112_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C4_N24112_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C4_N24112_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C4_N24112_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C12_N24114_O_3_C_6_io_in = {SBMux_C12_N24114_O_3_C_6_io_in_hi,SBMux_C12_N24114_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C12_N24114_O_3_C_6_io_config = configBlock_ioBundle_confOut[400:397]; // @[TileFull.scala 142:60]
  assign SBMux_C12_N24114_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C12_N24114_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C12_N24114_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C12_N24114_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C20_N24116_O_3_C_6_io_in = {SBMux_C20_N24116_O_3_C_6_io_in_hi,SBMux_C20_N24116_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C20_N24116_O_3_C_6_io_config = configBlock_ioBundle_confOut[404:401]; // @[TileFull.scala 142:60]
  assign SBMux_C20_N24116_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C20_N24116_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C20_N24116_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C20_N24116_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C28_N24118_O_3_C_6_io_in = {SBMux_C28_N24118_O_3_C_6_io_in_hi,SBMux_C28_N24118_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C28_N24118_O_3_C_6_io_config = configBlock_ioBundle_confOut[408:405]; // @[TileFull.scala 142:60]
  assign SBMux_C28_N24118_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C28_N24118_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C28_N24118_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C28_N24118_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C36_N24120_O_3_C_6_io_in = {SBMux_C36_N24120_O_3_C_6_io_in_hi,SBMux_C36_N24120_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C36_N24120_O_3_C_6_io_config = configBlock_ioBundle_confOut[412:409]; // @[TileFull.scala 142:60]
  assign SBMux_C36_N24120_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C36_N24120_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C36_N24120_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C36_N24120_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C44_N24122_O_4_C_5_io_in = {SBMux_C44_N24122_O_4_C_5_io_in_hi,SBMux_C44_N24122_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C44_N24122_O_4_C_5_io_config = configBlock_ioBundle_confOut[416:413]; // @[TileFull.scala 142:60]
  assign SBMux_C44_N24122_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C44_N24122_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C44_N24122_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C44_N24122_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C52_N24124_O_4_C_5_io_in = {SBMux_C52_N24124_O_4_C_5_io_in_hi,SBMux_C44_N24122_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C52_N24124_O_4_C_5_io_config = configBlock_ioBundle_confOut[420:417]; // @[TileFull.scala 142:60]
  assign SBMux_C52_N24124_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C52_N24124_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C52_N24124_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C52_N24124_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C60_N24126_O_4_C_5_io_in = {SBMux_C60_N24126_O_4_C_5_io_in_hi,SBMux_C60_N24126_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C60_N24126_O_4_C_5_io_config = configBlock_ioBundle_confOut[424:421]; // @[TileFull.scala 142:60]
  assign SBMux_C60_N24126_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C60_N24126_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C60_N24126_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C60_N24126_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C68_N24128_O_3_C_5_io_in = {SBMux_C68_N24128_O_3_C_5_io_in_hi,SBMux_C68_N24128_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C68_N24128_O_3_C_5_io_config = configBlock_ioBundle_confOut[428:425]; // @[TileFull.scala 142:60]
  assign SBMux_C68_N24128_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C68_N24128_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C68_N24128_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C68_N24128_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C76_N24130_O_0_C_4_io_in = {SBMux_C76_N24130_O_0_C_4_io_in_hi,SBMux_C76_N24130_O_0_C_4_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C76_N24130_O_0_C_4_io_config = configBlock_ioBundle_confOut[431:429]; // @[TileFull.scala 142:60]
  assign SBMux_C76_N24130_O_0_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C76_N24130_O_0_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C76_N24130_O_0_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C76_N24130_O_0_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C5_N27119_O_4_C_6_io_in = {SBMux_C5_N27119_O_4_C_6_io_in_hi,SBMux_C5_N27119_O_4_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C5_N27119_O_4_C_6_io_config = configBlock_ioBundle_confOut[435:432]; // @[TileFull.scala 142:60]
  assign SBMux_C5_N27119_O_4_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C5_N27119_O_4_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C5_N27119_O_4_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C5_N27119_O_4_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C13_N27127_O_3_C_6_io_in = {SBMux_C13_N27127_O_3_C_6_io_in_hi,SBMux_C13_N27127_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C13_N27127_O_3_C_6_io_config = configBlock_ioBundle_confOut[439:436]; // @[TileFull.scala 142:60]
  assign SBMux_C13_N27127_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C13_N27127_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C13_N27127_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C13_N27127_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C21_N27135_O_3_C_6_io_in = {SBMux_C21_N27135_O_3_C_6_io_in_hi,SBMux_C21_N27135_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C21_N27135_O_3_C_6_io_config = configBlock_ioBundle_confOut[443:440]; // @[TileFull.scala 142:60]
  assign SBMux_C21_N27135_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C21_N27135_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C21_N27135_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C21_N27135_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C29_N27143_O_3_C_5_io_in = {SBMux_C29_N27143_O_3_C_5_io_in_hi,SBMux_C29_N27143_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C29_N27143_O_3_C_5_io_config = configBlock_ioBundle_confOut[447:444]; // @[TileFull.scala 142:60]
  assign SBMux_C29_N27143_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C29_N27143_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C29_N27143_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C29_N27143_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C37_N27151_O_3_C_5_io_in = {SBMux_C37_N27151_O_3_C_5_io_in_hi,SBMux_C37_N27151_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C37_N27151_O_3_C_5_io_config = configBlock_ioBundle_confOut[451:448]; // @[TileFull.scala 142:60]
  assign SBMux_C37_N27151_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C37_N27151_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C37_N27151_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C37_N27151_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C45_N27159_O_4_C_5_io_in = {SBMux_C45_N27159_O_4_C_5_io_in_hi,SBMux_C45_N27159_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C45_N27159_O_4_C_5_io_config = configBlock_ioBundle_confOut[455:452]; // @[TileFull.scala 142:60]
  assign SBMux_C45_N27159_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C45_N27159_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C45_N27159_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C45_N27159_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C53_N27167_O_4_C_5_io_in = {SBMux_C53_N27167_O_4_C_5_io_in_hi,SBMux_C45_N27159_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C53_N27167_O_4_C_5_io_config = configBlock_ioBundle_confOut[459:456]; // @[TileFull.scala 142:60]
  assign SBMux_C53_N27167_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C53_N27167_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C53_N27167_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C53_N27167_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C61_N27175_O_4_C_5_io_in = {SBMux_C61_N27175_O_4_C_5_io_in_hi,SBMux_C61_N27175_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C61_N27175_O_4_C_5_io_config = configBlock_ioBundle_confOut[463:460]; // @[TileFull.scala 142:60]
  assign SBMux_C61_N27175_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C61_N27175_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C61_N27175_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C61_N27175_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C69_N27183_O_4_C_5_io_in = {SBMux_C69_N27183_O_4_C_5_io_in_hi,SBMux_C61_N27175_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C69_N27183_O_4_C_5_io_config = configBlock_ioBundle_confOut[467:464]; // @[TileFull.scala 142:60]
  assign SBMux_C69_N27183_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C69_N27183_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C69_N27183_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C69_N27183_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C77_N27215_O_3_C_5_io_in = {SBMux_C77_N27215_O_3_C_5_io_in_hi,SBMux_C77_N27215_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C77_N27215_O_3_C_5_io_config = configBlock_ioBundle_confOut[471:468]; // @[TileFull.scala 142:60]
  assign SBMux_C77_N27215_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C77_N27215_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C77_N27215_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C77_N27215_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C4_N27238_O_4_C_7_io_in = {SBMux_C4_N27238_O_4_C_7_io_in_hi,SBMux_C4_N27238_O_4_C_7_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C4_N27238_O_4_C_7_io_config = configBlock_ioBundle_confOut[475:472]; // @[TileFull.scala 142:60]
  assign SBMux_C4_N27238_O_4_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C4_N27238_O_4_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C4_N27238_O_4_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C4_N27238_O_4_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C12_N27240_O_3_C_6_io_in = {SBMux_C12_N27240_O_3_C_6_io_in_hi,SBMux_C12_N27240_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C12_N27240_O_3_C_6_io_config = configBlock_ioBundle_confOut[479:476]; // @[TileFull.scala 142:60]
  assign SBMux_C12_N27240_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C12_N27240_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C12_N27240_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C12_N27240_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C20_N27242_O_3_C_6_io_in = {SBMux_C20_N27242_O_3_C_6_io_in_hi,SBMux_C20_N27242_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C20_N27242_O_3_C_6_io_config = configBlock_ioBundle_confOut[483:480]; // @[TileFull.scala 142:60]
  assign SBMux_C20_N27242_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C20_N27242_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C20_N27242_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C20_N27242_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C28_N27244_O_3_C_5_io_in = {SBMux_C28_N27244_O_3_C_5_io_in_hi,SBMux_C28_N27244_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C28_N27244_O_3_C_5_io_config = configBlock_ioBundle_confOut[487:484]; // @[TileFull.scala 142:60]
  assign SBMux_C28_N27244_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C28_N27244_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C28_N27244_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C28_N27244_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C36_N27246_O_3_C_5_io_in = {SBMux_C36_N27246_O_3_C_5_io_in_hi,SBMux_C36_N27246_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C36_N27246_O_3_C_5_io_config = configBlock_ioBundle_confOut[491:488]; // @[TileFull.scala 142:60]
  assign SBMux_C36_N27246_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C36_N27246_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C36_N27246_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C36_N27246_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C44_N27248_O_4_C_5_io_in = {SBMux_C44_N27248_O_4_C_5_io_in_hi,SBMux_C44_N27248_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C44_N27248_O_4_C_5_io_config = configBlock_ioBundle_confOut[495:492]; // @[TileFull.scala 142:60]
  assign SBMux_C44_N27248_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C44_N27248_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C44_N27248_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C44_N27248_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C52_N27250_O_4_C_5_io_in = {SBMux_C52_N27250_O_4_C_5_io_in_hi,SBMux_C44_N27248_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C52_N27250_O_4_C_5_io_config = configBlock_ioBundle_confOut[499:496]; // @[TileFull.scala 142:60]
  assign SBMux_C52_N27250_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C52_N27250_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C52_N27250_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C52_N27250_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C60_N27252_O_4_C_6_io_in = {SBMux_C60_N27252_O_4_C_6_io_in_hi,SBMux_C60_N27252_O_4_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C60_N27252_O_4_C_6_io_config = configBlock_ioBundle_confOut[503:500]; // @[TileFull.scala 142:60]
  assign SBMux_C60_N27252_O_4_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C60_N27252_O_4_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C60_N27252_O_4_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C60_N27252_O_4_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C68_N27254_O_4_C_6_io_in = {SBMux_C68_N27254_O_4_C_6_io_in_hi,SBMux_C68_N27254_O_4_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C68_N27254_O_4_C_6_io_config = configBlock_ioBundle_confOut[507:504]; // @[TileFull.scala 142:60]
  assign SBMux_C68_N27254_O_4_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C68_N27254_O_4_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C68_N27254_O_4_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C68_N27254_O_4_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C76_N27256_O_3_C_7_io_in = {SBMux_C76_N27256_O_3_C_7_io_in_hi,SBMux_C76_N27256_O_3_C_7_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C76_N27256_O_3_C_7_io_config = configBlock_ioBundle_confOut[511:508]; // @[TileFull.scala 142:60]
  assign SBMux_C76_N27256_O_3_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C76_N27256_O_3_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C76_N27256_O_3_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C76_N27256_O_3_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
endmodule
