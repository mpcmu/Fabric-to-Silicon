/afs/ece.cmu.edu/project/km_group/.vol9/asap7/asap7sc7p5t_28/LEF/scaled/asap7sc7p5t_28_SRAM_4x_220121a.lef