module IOBlock(
  input         IPIN_0,
  input         IPIN_2,
  input         IPIN_4,
  input         IPIN_6,
  input         IPIN_8,
  input         IPIN_10,
  input         IPIN_12,
  input         IPIN_14,
  input         IPIN_16,
  input         IPIN_18,
  input         IPIN_20,
  input         IPIN_22,
  input         IPIN_24,
  input         IPIN_26,
  input         IPIN_28,
  input         IPIN_30,
  input         IPIN_32,
  input         IPIN_34,
  input         IPIN_36,
  input         IPIN_38,
  input         IPIN_40,
  input         IPIN_42,
  input         IPIN_44,
  input         IPIN_46,
  input         IPIN_48,
  input         IPIN_50,
  input         IPIN_52,
  input         IPIN_54,
  input         IPIN_56,
  input         IPIN_58,
  input         IPIN_60,
  input         IPIN_62,
  output        OPIN_1,
  output        OPIN_3,
  output        OPIN_5,
  output        OPIN_7,
  output        OPIN_9,
  output        OPIN_11,
  output        OPIN_13,
  output        OPIN_15,
  output        OPIN_17,
  output        OPIN_19,
  output        OPIN_21,
  output        OPIN_23,
  output        OPIN_25,
  output        OPIN_27,
  output        OPIN_29,
  output        OPIN_31,
  output        OPIN_33,
  output        OPIN_35,
  output        OPIN_37,
  output        OPIN_39,
  output        OPIN_41,
  output        OPIN_43,
  output        OPIN_45,
  output        OPIN_47,
  output        OPIN_49,
  output        OPIN_51,
  output        OPIN_53,
  output        OPIN_55,
  output        OPIN_57,
  output        OPIN_59,
  output        OPIN_61,
  output        OPIN_63,
  input         clock,
  input         reset,
  input  [31:0] ioPad_i,
  output [31:0] ioPad_o,
  input  [15:0] configBits,
  input         loopBreak,
  input         gndLBouts
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] padOutReg_lo_lo = {IPIN_14,IPIN_12,IPIN_10,IPIN_8,IPIN_6,IPIN_4,IPIN_2,IPIN_0}; // @[IOBlock.scala 31:60]
  wire [15:0] padOutReg_lo = {IPIN_30,IPIN_28,IPIN_26,IPIN_24,IPIN_22,IPIN_20,IPIN_18,IPIN_16,padOutReg_lo_lo}; // @[IOBlock.scala 31:60]
  wire [7:0] padOutReg_hi_lo = {IPIN_46,IPIN_44,IPIN_42,IPIN_40,IPIN_38,IPIN_36,IPIN_34,IPIN_32}; // @[IOBlock.scala 31:60]
  wire [31:0] _padOutReg_T = {IPIN_62,IPIN_60,IPIN_58,IPIN_56,IPIN_54,IPIN_52,IPIN_50,IPIN_48,padOutReg_hi_lo,
    padOutReg_lo}; // @[IOBlock.scala 31:60]
  reg [31:0] padOutReg; // @[Reg.scala 28:20]
  wire [31:0] padOut = loopBreak ? padOutReg : _padOutReg_T; // @[IOBlock.scala 32:21]
  reg [31:0] padInReg; // @[IOBlock.scala 36:27]
  reg [31:0] padInReg_r; // @[Reg.scala 28:20]
  wire [31:0] _padIn_T = loopBreak ? padInReg : ioPad_i; // @[IOBlock.scala 38:40]
  wire [31:0] padIn = gndLBouts ? 32'h0 : _padIn_T; // @[IOBlock.scala 38:20]
  assign OPIN_1 = padIn[0]; // @[IOBlock.scala 45:28]
  assign OPIN_3 = padIn[1]; // @[IOBlock.scala 45:28]
  assign OPIN_5 = padIn[2]; // @[IOBlock.scala 45:28]
  assign OPIN_7 = padIn[3]; // @[IOBlock.scala 45:28]
  assign OPIN_9 = padIn[4]; // @[IOBlock.scala 45:28]
  assign OPIN_11 = padIn[5]; // @[IOBlock.scala 45:28]
  assign OPIN_13 = padIn[6]; // @[IOBlock.scala 45:28]
  assign OPIN_15 = padIn[7]; // @[IOBlock.scala 45:28]
  assign OPIN_17 = padIn[8]; // @[IOBlock.scala 45:28]
  assign OPIN_19 = padIn[9]; // @[IOBlock.scala 45:28]
  assign OPIN_21 = padIn[10]; // @[IOBlock.scala 45:28]
  assign OPIN_23 = padIn[11]; // @[IOBlock.scala 45:28]
  assign OPIN_25 = padIn[12]; // @[IOBlock.scala 45:28]
  assign OPIN_27 = padIn[13]; // @[IOBlock.scala 45:28]
  assign OPIN_29 = padIn[14]; // @[IOBlock.scala 45:28]
  assign OPIN_31 = padIn[15]; // @[IOBlock.scala 45:28]
  assign OPIN_33 = padIn[16]; // @[IOBlock.scala 45:28]
  assign OPIN_35 = padIn[17]; // @[IOBlock.scala 45:28]
  assign OPIN_37 = padIn[18]; // @[IOBlock.scala 45:28]
  assign OPIN_39 = padIn[19]; // @[IOBlock.scala 45:28]
  assign OPIN_41 = padIn[20]; // @[IOBlock.scala 45:28]
  assign OPIN_43 = padIn[21]; // @[IOBlock.scala 45:28]
  assign OPIN_45 = padIn[22]; // @[IOBlock.scala 45:28]
  assign OPIN_47 = padIn[23]; // @[IOBlock.scala 45:28]
  assign OPIN_49 = padIn[24]; // @[IOBlock.scala 45:28]
  assign OPIN_51 = padIn[25]; // @[IOBlock.scala 45:28]
  assign OPIN_53 = padIn[26]; // @[IOBlock.scala 45:28]
  assign OPIN_55 = padIn[27]; // @[IOBlock.scala 45:28]
  assign OPIN_57 = padIn[28]; // @[IOBlock.scala 45:28]
  assign OPIN_59 = padIn[29]; // @[IOBlock.scala 45:28]
  assign OPIN_61 = padIn[30]; // @[IOBlock.scala 45:28]
  assign OPIN_63 = padIn[31]; // @[IOBlock.scala 45:28]
  assign ioPad_o = gndLBouts ? 32'h0 : padOut; // @[IOBlock.scala 33:23]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      padOutReg <= 32'h0; // @[Reg.scala 28:20]
    end else if (configBits[15]) begin // @[Reg.scala 29:18]
      padOutReg <= _padOutReg_T; // @[Reg.scala 29:22]
    end
    if (reset) begin // @[IOBlock.scala 36:27]
      padInReg <= 32'h0; // @[IOBlock.scala 36:27]
    end else begin
      padInReg <= padInReg_r; // @[IOBlock.scala 37:14]
    end
    if (reset) begin // @[Reg.scala 28:20]
      padInReg_r <= 32'h0; // @[Reg.scala 28:20]
    end else if (configBits[15]) begin // @[Reg.scala 29:18]
      padInReg_r <= ioPad_i; // @[Reg.scala 29:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  padOutReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  padInReg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  padInReg_r = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ScanConf_Tile_11_3_iotile(
  input          clock,
  output [423:0] ioBundle_confOut,
  input  [7:0]   ioBundle_scan_in,
  input          ioBundle_scan_en,
  output [7:0]   ioBundle_scan_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
`endif // RANDOMIZE_REG_INIT
  reg  confReg_0; // @[ScanConf.scala 32:20]
  reg  confReg_1; // @[ScanConf.scala 32:20]
  reg  confReg_2; // @[ScanConf.scala 32:20]
  reg  confReg_3; // @[ScanConf.scala 32:20]
  reg  confReg_4; // @[ScanConf.scala 32:20]
  reg  confReg_5; // @[ScanConf.scala 32:20]
  reg  confReg_6; // @[ScanConf.scala 32:20]
  reg  confReg_7; // @[ScanConf.scala 32:20]
  reg  confReg_8; // @[ScanConf.scala 32:20]
  reg  confReg_9; // @[ScanConf.scala 32:20]
  reg  confReg_10; // @[ScanConf.scala 32:20]
  reg  confReg_11; // @[ScanConf.scala 32:20]
  reg  confReg_12; // @[ScanConf.scala 32:20]
  reg  confReg_13; // @[ScanConf.scala 32:20]
  reg  confReg_14; // @[ScanConf.scala 32:20]
  reg  confReg_15; // @[ScanConf.scala 32:20]
  reg  confReg_16; // @[ScanConf.scala 32:20]
  reg  confReg_17; // @[ScanConf.scala 32:20]
  reg  confReg_18; // @[ScanConf.scala 32:20]
  reg  confReg_19; // @[ScanConf.scala 32:20]
  reg  confReg_20; // @[ScanConf.scala 32:20]
  reg  confReg_21; // @[ScanConf.scala 32:20]
  reg  confReg_22; // @[ScanConf.scala 32:20]
  reg  confReg_23; // @[ScanConf.scala 32:20]
  reg  confReg_24; // @[ScanConf.scala 32:20]
  reg  confReg_25; // @[ScanConf.scala 32:20]
  reg  confReg_26; // @[ScanConf.scala 32:20]
  reg  confReg_27; // @[ScanConf.scala 32:20]
  reg  confReg_28; // @[ScanConf.scala 32:20]
  reg  confReg_29; // @[ScanConf.scala 32:20]
  reg  confReg_30; // @[ScanConf.scala 32:20]
  reg  confReg_31; // @[ScanConf.scala 32:20]
  reg  confReg_32; // @[ScanConf.scala 32:20]
  reg  confReg_33; // @[ScanConf.scala 32:20]
  reg  confReg_34; // @[ScanConf.scala 32:20]
  reg  confReg_35; // @[ScanConf.scala 32:20]
  reg  confReg_36; // @[ScanConf.scala 32:20]
  reg  confReg_37; // @[ScanConf.scala 32:20]
  reg  confReg_38; // @[ScanConf.scala 32:20]
  reg  confReg_39; // @[ScanConf.scala 32:20]
  reg  confReg_40; // @[ScanConf.scala 32:20]
  reg  confReg_41; // @[ScanConf.scala 32:20]
  reg  confReg_42; // @[ScanConf.scala 32:20]
  reg  confReg_43; // @[ScanConf.scala 32:20]
  reg  confReg_44; // @[ScanConf.scala 32:20]
  reg  confReg_45; // @[ScanConf.scala 32:20]
  reg  confReg_46; // @[ScanConf.scala 32:20]
  reg  confReg_47; // @[ScanConf.scala 32:20]
  reg  confReg_48; // @[ScanConf.scala 32:20]
  reg  confReg_49; // @[ScanConf.scala 32:20]
  reg  confReg_50; // @[ScanConf.scala 32:20]
  reg  confReg_51; // @[ScanConf.scala 32:20]
  reg  confReg_52; // @[ScanConf.scala 32:20]
  reg  confReg_53; // @[ScanConf.scala 32:20]
  reg  confReg_54; // @[ScanConf.scala 32:20]
  reg  confReg_55; // @[ScanConf.scala 32:20]
  reg  confReg_56; // @[ScanConf.scala 32:20]
  reg  confReg_57; // @[ScanConf.scala 32:20]
  reg  confReg_58; // @[ScanConf.scala 32:20]
  reg  confReg_59; // @[ScanConf.scala 32:20]
  reg  confReg_60; // @[ScanConf.scala 32:20]
  reg  confReg_61; // @[ScanConf.scala 32:20]
  reg  confReg_62; // @[ScanConf.scala 32:20]
  reg  confReg_63; // @[ScanConf.scala 32:20]
  reg  confReg_64; // @[ScanConf.scala 32:20]
  reg  confReg_65; // @[ScanConf.scala 32:20]
  reg  confReg_66; // @[ScanConf.scala 32:20]
  reg  confReg_67; // @[ScanConf.scala 32:20]
  reg  confReg_68; // @[ScanConf.scala 32:20]
  reg  confReg_69; // @[ScanConf.scala 32:20]
  reg  confReg_70; // @[ScanConf.scala 32:20]
  reg  confReg_71; // @[ScanConf.scala 32:20]
  reg  confReg_72; // @[ScanConf.scala 32:20]
  reg  confReg_73; // @[ScanConf.scala 32:20]
  reg  confReg_74; // @[ScanConf.scala 32:20]
  reg  confReg_75; // @[ScanConf.scala 32:20]
  reg  confReg_76; // @[ScanConf.scala 32:20]
  reg  confReg_77; // @[ScanConf.scala 32:20]
  reg  confReg_78; // @[ScanConf.scala 32:20]
  reg  confReg_79; // @[ScanConf.scala 32:20]
  reg  confReg_80; // @[ScanConf.scala 32:20]
  reg  confReg_81; // @[ScanConf.scala 32:20]
  reg  confReg_82; // @[ScanConf.scala 32:20]
  reg  confReg_83; // @[ScanConf.scala 32:20]
  reg  confReg_84; // @[ScanConf.scala 32:20]
  reg  confReg_85; // @[ScanConf.scala 32:20]
  reg  confReg_86; // @[ScanConf.scala 32:20]
  reg  confReg_87; // @[ScanConf.scala 32:20]
  reg  confReg_88; // @[ScanConf.scala 32:20]
  reg  confReg_89; // @[ScanConf.scala 32:20]
  reg  confReg_90; // @[ScanConf.scala 32:20]
  reg  confReg_91; // @[ScanConf.scala 32:20]
  reg  confReg_92; // @[ScanConf.scala 32:20]
  reg  confReg_93; // @[ScanConf.scala 32:20]
  reg  confReg_94; // @[ScanConf.scala 32:20]
  reg  confReg_95; // @[ScanConf.scala 32:20]
  reg  confReg_96; // @[ScanConf.scala 32:20]
  reg  confReg_97; // @[ScanConf.scala 32:20]
  reg  confReg_98; // @[ScanConf.scala 32:20]
  reg  confReg_99; // @[ScanConf.scala 32:20]
  reg  confReg_100; // @[ScanConf.scala 32:20]
  reg  confReg_101; // @[ScanConf.scala 32:20]
  reg  confReg_102; // @[ScanConf.scala 32:20]
  reg  confReg_103; // @[ScanConf.scala 32:20]
  reg  confReg_104; // @[ScanConf.scala 32:20]
  reg  confReg_105; // @[ScanConf.scala 32:20]
  reg  confReg_106; // @[ScanConf.scala 32:20]
  reg  confReg_107; // @[ScanConf.scala 32:20]
  reg  confReg_108; // @[ScanConf.scala 32:20]
  reg  confReg_109; // @[ScanConf.scala 32:20]
  reg  confReg_110; // @[ScanConf.scala 32:20]
  reg  confReg_111; // @[ScanConf.scala 32:20]
  reg  confReg_112; // @[ScanConf.scala 32:20]
  reg  confReg_113; // @[ScanConf.scala 32:20]
  reg  confReg_114; // @[ScanConf.scala 32:20]
  reg  confReg_115; // @[ScanConf.scala 32:20]
  reg  confReg_116; // @[ScanConf.scala 32:20]
  reg  confReg_117; // @[ScanConf.scala 32:20]
  reg  confReg_118; // @[ScanConf.scala 32:20]
  reg  confReg_119; // @[ScanConf.scala 32:20]
  reg  confReg_120; // @[ScanConf.scala 32:20]
  reg  confReg_121; // @[ScanConf.scala 32:20]
  reg  confReg_122; // @[ScanConf.scala 32:20]
  reg  confReg_123; // @[ScanConf.scala 32:20]
  reg  confReg_124; // @[ScanConf.scala 32:20]
  reg  confReg_125; // @[ScanConf.scala 32:20]
  reg  confReg_126; // @[ScanConf.scala 32:20]
  reg  confReg_127; // @[ScanConf.scala 32:20]
  reg  confReg_128; // @[ScanConf.scala 32:20]
  reg  confReg_129; // @[ScanConf.scala 32:20]
  reg  confReg_130; // @[ScanConf.scala 32:20]
  reg  confReg_131; // @[ScanConf.scala 32:20]
  reg  confReg_132; // @[ScanConf.scala 32:20]
  reg  confReg_133; // @[ScanConf.scala 32:20]
  reg  confReg_134; // @[ScanConf.scala 32:20]
  reg  confReg_135; // @[ScanConf.scala 32:20]
  reg  confReg_136; // @[ScanConf.scala 32:20]
  reg  confReg_137; // @[ScanConf.scala 32:20]
  reg  confReg_138; // @[ScanConf.scala 32:20]
  reg  confReg_139; // @[ScanConf.scala 32:20]
  reg  confReg_140; // @[ScanConf.scala 32:20]
  reg  confReg_141; // @[ScanConf.scala 32:20]
  reg  confReg_142; // @[ScanConf.scala 32:20]
  reg  confReg_143; // @[ScanConf.scala 32:20]
  reg  confReg_144; // @[ScanConf.scala 32:20]
  reg  confReg_145; // @[ScanConf.scala 32:20]
  reg  confReg_146; // @[ScanConf.scala 32:20]
  reg  confReg_147; // @[ScanConf.scala 32:20]
  reg  confReg_148; // @[ScanConf.scala 32:20]
  reg  confReg_149; // @[ScanConf.scala 32:20]
  reg  confReg_150; // @[ScanConf.scala 32:20]
  reg  confReg_151; // @[ScanConf.scala 32:20]
  reg  confReg_152; // @[ScanConf.scala 32:20]
  reg  confReg_153; // @[ScanConf.scala 32:20]
  reg  confReg_154; // @[ScanConf.scala 32:20]
  reg  confReg_155; // @[ScanConf.scala 32:20]
  reg  confReg_156; // @[ScanConf.scala 32:20]
  reg  confReg_157; // @[ScanConf.scala 32:20]
  reg  confReg_158; // @[ScanConf.scala 32:20]
  reg  confReg_159; // @[ScanConf.scala 32:20]
  reg  confReg_160; // @[ScanConf.scala 32:20]
  reg  confReg_161; // @[ScanConf.scala 32:20]
  reg  confReg_162; // @[ScanConf.scala 32:20]
  reg  confReg_163; // @[ScanConf.scala 32:20]
  reg  confReg_164; // @[ScanConf.scala 32:20]
  reg  confReg_165; // @[ScanConf.scala 32:20]
  reg  confReg_166; // @[ScanConf.scala 32:20]
  reg  confReg_167; // @[ScanConf.scala 32:20]
  reg  confReg_168; // @[ScanConf.scala 32:20]
  reg  confReg_169; // @[ScanConf.scala 32:20]
  reg  confReg_170; // @[ScanConf.scala 32:20]
  reg  confReg_171; // @[ScanConf.scala 32:20]
  reg  confReg_172; // @[ScanConf.scala 32:20]
  reg  confReg_173; // @[ScanConf.scala 32:20]
  reg  confReg_174; // @[ScanConf.scala 32:20]
  reg  confReg_175; // @[ScanConf.scala 32:20]
  reg  confReg_176; // @[ScanConf.scala 32:20]
  reg  confReg_177; // @[ScanConf.scala 32:20]
  reg  confReg_178; // @[ScanConf.scala 32:20]
  reg  confReg_179; // @[ScanConf.scala 32:20]
  reg  confReg_180; // @[ScanConf.scala 32:20]
  reg  confReg_181; // @[ScanConf.scala 32:20]
  reg  confReg_182; // @[ScanConf.scala 32:20]
  reg  confReg_183; // @[ScanConf.scala 32:20]
  reg  confReg_184; // @[ScanConf.scala 32:20]
  reg  confReg_185; // @[ScanConf.scala 32:20]
  reg  confReg_186; // @[ScanConf.scala 32:20]
  reg  confReg_187; // @[ScanConf.scala 32:20]
  reg  confReg_188; // @[ScanConf.scala 32:20]
  reg  confReg_189; // @[ScanConf.scala 32:20]
  reg  confReg_190; // @[ScanConf.scala 32:20]
  reg  confReg_191; // @[ScanConf.scala 32:20]
  reg  confReg_192; // @[ScanConf.scala 32:20]
  reg  confReg_193; // @[ScanConf.scala 32:20]
  reg  confReg_194; // @[ScanConf.scala 32:20]
  reg  confReg_195; // @[ScanConf.scala 32:20]
  reg  confReg_196; // @[ScanConf.scala 32:20]
  reg  confReg_197; // @[ScanConf.scala 32:20]
  reg  confReg_198; // @[ScanConf.scala 32:20]
  reg  confReg_199; // @[ScanConf.scala 32:20]
  reg  confReg_200; // @[ScanConf.scala 32:20]
  reg  confReg_201; // @[ScanConf.scala 32:20]
  reg  confReg_202; // @[ScanConf.scala 32:20]
  reg  confReg_203; // @[ScanConf.scala 32:20]
  reg  confReg_204; // @[ScanConf.scala 32:20]
  reg  confReg_205; // @[ScanConf.scala 32:20]
  reg  confReg_206; // @[ScanConf.scala 32:20]
  reg  confReg_207; // @[ScanConf.scala 32:20]
  reg  confReg_208; // @[ScanConf.scala 32:20]
  reg  confReg_209; // @[ScanConf.scala 32:20]
  reg  confReg_210; // @[ScanConf.scala 32:20]
  reg  confReg_211; // @[ScanConf.scala 32:20]
  reg  confReg_212; // @[ScanConf.scala 32:20]
  reg  confReg_213; // @[ScanConf.scala 32:20]
  reg  confReg_214; // @[ScanConf.scala 32:20]
  reg  confReg_215; // @[ScanConf.scala 32:20]
  reg  confReg_216; // @[ScanConf.scala 32:20]
  reg  confReg_217; // @[ScanConf.scala 32:20]
  reg  confReg_218; // @[ScanConf.scala 32:20]
  reg  confReg_219; // @[ScanConf.scala 32:20]
  reg  confReg_220; // @[ScanConf.scala 32:20]
  reg  confReg_221; // @[ScanConf.scala 32:20]
  reg  confReg_222; // @[ScanConf.scala 32:20]
  reg  confReg_223; // @[ScanConf.scala 32:20]
  reg  confReg_224; // @[ScanConf.scala 32:20]
  reg  confReg_225; // @[ScanConf.scala 32:20]
  reg  confReg_226; // @[ScanConf.scala 32:20]
  reg  confReg_227; // @[ScanConf.scala 32:20]
  reg  confReg_228; // @[ScanConf.scala 32:20]
  reg  confReg_229; // @[ScanConf.scala 32:20]
  reg  confReg_230; // @[ScanConf.scala 32:20]
  reg  confReg_231; // @[ScanConf.scala 32:20]
  reg  confReg_232; // @[ScanConf.scala 32:20]
  reg  confReg_233; // @[ScanConf.scala 32:20]
  reg  confReg_234; // @[ScanConf.scala 32:20]
  reg  confReg_235; // @[ScanConf.scala 32:20]
  reg  confReg_236; // @[ScanConf.scala 32:20]
  reg  confReg_237; // @[ScanConf.scala 32:20]
  reg  confReg_238; // @[ScanConf.scala 32:20]
  reg  confReg_239; // @[ScanConf.scala 32:20]
  reg  confReg_240; // @[ScanConf.scala 32:20]
  reg  confReg_241; // @[ScanConf.scala 32:20]
  reg  confReg_242; // @[ScanConf.scala 32:20]
  reg  confReg_243; // @[ScanConf.scala 32:20]
  reg  confReg_244; // @[ScanConf.scala 32:20]
  reg  confReg_245; // @[ScanConf.scala 32:20]
  reg  confReg_246; // @[ScanConf.scala 32:20]
  reg  confReg_247; // @[ScanConf.scala 32:20]
  reg  confReg_248; // @[ScanConf.scala 32:20]
  reg  confReg_249; // @[ScanConf.scala 32:20]
  reg  confReg_250; // @[ScanConf.scala 32:20]
  reg  confReg_251; // @[ScanConf.scala 32:20]
  reg  confReg_252; // @[ScanConf.scala 32:20]
  reg  confReg_253; // @[ScanConf.scala 32:20]
  reg  confReg_254; // @[ScanConf.scala 32:20]
  reg  confReg_255; // @[ScanConf.scala 32:20]
  reg  confReg_256; // @[ScanConf.scala 32:20]
  reg  confReg_257; // @[ScanConf.scala 32:20]
  reg  confReg_258; // @[ScanConf.scala 32:20]
  reg  confReg_259; // @[ScanConf.scala 32:20]
  reg  confReg_260; // @[ScanConf.scala 32:20]
  reg  confReg_261; // @[ScanConf.scala 32:20]
  reg  confReg_262; // @[ScanConf.scala 32:20]
  reg  confReg_263; // @[ScanConf.scala 32:20]
  reg  confReg_264; // @[ScanConf.scala 32:20]
  reg  confReg_265; // @[ScanConf.scala 32:20]
  reg  confReg_266; // @[ScanConf.scala 32:20]
  reg  confReg_267; // @[ScanConf.scala 32:20]
  reg  confReg_268; // @[ScanConf.scala 32:20]
  reg  confReg_269; // @[ScanConf.scala 32:20]
  reg  confReg_270; // @[ScanConf.scala 32:20]
  reg  confReg_271; // @[ScanConf.scala 32:20]
  reg  confReg_272; // @[ScanConf.scala 32:20]
  reg  confReg_273; // @[ScanConf.scala 32:20]
  reg  confReg_274; // @[ScanConf.scala 32:20]
  reg  confReg_275; // @[ScanConf.scala 32:20]
  reg  confReg_276; // @[ScanConf.scala 32:20]
  reg  confReg_277; // @[ScanConf.scala 32:20]
  reg  confReg_278; // @[ScanConf.scala 32:20]
  reg  confReg_279; // @[ScanConf.scala 32:20]
  reg  confReg_280; // @[ScanConf.scala 32:20]
  reg  confReg_281; // @[ScanConf.scala 32:20]
  reg  confReg_282; // @[ScanConf.scala 32:20]
  reg  confReg_283; // @[ScanConf.scala 32:20]
  reg  confReg_284; // @[ScanConf.scala 32:20]
  reg  confReg_285; // @[ScanConf.scala 32:20]
  reg  confReg_286; // @[ScanConf.scala 32:20]
  reg  confReg_287; // @[ScanConf.scala 32:20]
  reg  confReg_288; // @[ScanConf.scala 32:20]
  reg  confReg_289; // @[ScanConf.scala 32:20]
  reg  confReg_290; // @[ScanConf.scala 32:20]
  reg  confReg_291; // @[ScanConf.scala 32:20]
  reg  confReg_292; // @[ScanConf.scala 32:20]
  reg  confReg_293; // @[ScanConf.scala 32:20]
  reg  confReg_294; // @[ScanConf.scala 32:20]
  reg  confReg_295; // @[ScanConf.scala 32:20]
  reg  confReg_296; // @[ScanConf.scala 32:20]
  reg  confReg_297; // @[ScanConf.scala 32:20]
  reg  confReg_298; // @[ScanConf.scala 32:20]
  reg  confReg_299; // @[ScanConf.scala 32:20]
  reg  confReg_300; // @[ScanConf.scala 32:20]
  reg  confReg_301; // @[ScanConf.scala 32:20]
  reg  confReg_302; // @[ScanConf.scala 32:20]
  reg  confReg_303; // @[ScanConf.scala 32:20]
  reg  confReg_304; // @[ScanConf.scala 32:20]
  reg  confReg_305; // @[ScanConf.scala 32:20]
  reg  confReg_306; // @[ScanConf.scala 32:20]
  reg  confReg_307; // @[ScanConf.scala 32:20]
  reg  confReg_308; // @[ScanConf.scala 32:20]
  reg  confReg_309; // @[ScanConf.scala 32:20]
  reg  confReg_310; // @[ScanConf.scala 32:20]
  reg  confReg_311; // @[ScanConf.scala 32:20]
  reg  confReg_312; // @[ScanConf.scala 32:20]
  reg  confReg_313; // @[ScanConf.scala 32:20]
  reg  confReg_314; // @[ScanConf.scala 32:20]
  reg  confReg_315; // @[ScanConf.scala 32:20]
  reg  confReg_316; // @[ScanConf.scala 32:20]
  reg  confReg_317; // @[ScanConf.scala 32:20]
  reg  confReg_318; // @[ScanConf.scala 32:20]
  reg  confReg_319; // @[ScanConf.scala 32:20]
  reg  confReg_320; // @[ScanConf.scala 32:20]
  reg  confReg_321; // @[ScanConf.scala 32:20]
  reg  confReg_322; // @[ScanConf.scala 32:20]
  reg  confReg_323; // @[ScanConf.scala 32:20]
  reg  confReg_324; // @[ScanConf.scala 32:20]
  reg  confReg_325; // @[ScanConf.scala 32:20]
  reg  confReg_326; // @[ScanConf.scala 32:20]
  reg  confReg_327; // @[ScanConf.scala 32:20]
  reg  confReg_328; // @[ScanConf.scala 32:20]
  reg  confReg_329; // @[ScanConf.scala 32:20]
  reg  confReg_330; // @[ScanConf.scala 32:20]
  reg  confReg_331; // @[ScanConf.scala 32:20]
  reg  confReg_332; // @[ScanConf.scala 32:20]
  reg  confReg_333; // @[ScanConf.scala 32:20]
  reg  confReg_334; // @[ScanConf.scala 32:20]
  reg  confReg_335; // @[ScanConf.scala 32:20]
  reg  confReg_336; // @[ScanConf.scala 32:20]
  reg  confReg_337; // @[ScanConf.scala 32:20]
  reg  confReg_338; // @[ScanConf.scala 32:20]
  reg  confReg_339; // @[ScanConf.scala 32:20]
  reg  confReg_340; // @[ScanConf.scala 32:20]
  reg  confReg_341; // @[ScanConf.scala 32:20]
  reg  confReg_342; // @[ScanConf.scala 32:20]
  reg  confReg_343; // @[ScanConf.scala 32:20]
  reg  confReg_344; // @[ScanConf.scala 32:20]
  reg  confReg_345; // @[ScanConf.scala 32:20]
  reg  confReg_346; // @[ScanConf.scala 32:20]
  reg  confReg_347; // @[ScanConf.scala 32:20]
  reg  confReg_348; // @[ScanConf.scala 32:20]
  reg  confReg_349; // @[ScanConf.scala 32:20]
  reg  confReg_350; // @[ScanConf.scala 32:20]
  reg  confReg_351; // @[ScanConf.scala 32:20]
  reg  confReg_352; // @[ScanConf.scala 32:20]
  reg  confReg_353; // @[ScanConf.scala 32:20]
  reg  confReg_354; // @[ScanConf.scala 32:20]
  reg  confReg_355; // @[ScanConf.scala 32:20]
  reg  confReg_356; // @[ScanConf.scala 32:20]
  reg  confReg_357; // @[ScanConf.scala 32:20]
  reg  confReg_358; // @[ScanConf.scala 32:20]
  reg  confReg_359; // @[ScanConf.scala 32:20]
  reg  confReg_360; // @[ScanConf.scala 32:20]
  reg  confReg_361; // @[ScanConf.scala 32:20]
  reg  confReg_362; // @[ScanConf.scala 32:20]
  reg  confReg_363; // @[ScanConf.scala 32:20]
  reg  confReg_364; // @[ScanConf.scala 32:20]
  reg  confReg_365; // @[ScanConf.scala 32:20]
  reg  confReg_366; // @[ScanConf.scala 32:20]
  reg  confReg_367; // @[ScanConf.scala 32:20]
  reg  confReg_368; // @[ScanConf.scala 32:20]
  reg  confReg_369; // @[ScanConf.scala 32:20]
  reg  confReg_370; // @[ScanConf.scala 32:20]
  reg  confReg_371; // @[ScanConf.scala 32:20]
  reg  confReg_372; // @[ScanConf.scala 32:20]
  reg  confReg_373; // @[ScanConf.scala 32:20]
  reg  confReg_374; // @[ScanConf.scala 32:20]
  reg  confReg_375; // @[ScanConf.scala 32:20]
  reg  confReg_376; // @[ScanConf.scala 32:20]
  reg  confReg_377; // @[ScanConf.scala 32:20]
  reg  confReg_378; // @[ScanConf.scala 32:20]
  reg  confReg_379; // @[ScanConf.scala 32:20]
  reg  confReg_380; // @[ScanConf.scala 32:20]
  reg  confReg_381; // @[ScanConf.scala 32:20]
  reg  confReg_382; // @[ScanConf.scala 32:20]
  reg  confReg_383; // @[ScanConf.scala 32:20]
  reg  confReg_384; // @[ScanConf.scala 32:20]
  reg  confReg_385; // @[ScanConf.scala 32:20]
  reg  confReg_386; // @[ScanConf.scala 32:20]
  reg  confReg_387; // @[ScanConf.scala 32:20]
  reg  confReg_388; // @[ScanConf.scala 32:20]
  reg  confReg_389; // @[ScanConf.scala 32:20]
  reg  confReg_390; // @[ScanConf.scala 32:20]
  reg  confReg_391; // @[ScanConf.scala 32:20]
  reg  confReg_392; // @[ScanConf.scala 32:20]
  reg  confReg_393; // @[ScanConf.scala 32:20]
  reg  confReg_394; // @[ScanConf.scala 32:20]
  reg  confReg_395; // @[ScanConf.scala 32:20]
  reg  confReg_396; // @[ScanConf.scala 32:20]
  reg  confReg_397; // @[ScanConf.scala 32:20]
  reg  confReg_398; // @[ScanConf.scala 32:20]
  reg  confReg_399; // @[ScanConf.scala 32:20]
  reg  confReg_400; // @[ScanConf.scala 32:20]
  reg  confReg_401; // @[ScanConf.scala 32:20]
  reg  confReg_402; // @[ScanConf.scala 32:20]
  reg  confReg_403; // @[ScanConf.scala 32:20]
  reg  confReg_404; // @[ScanConf.scala 32:20]
  reg  confReg_405; // @[ScanConf.scala 32:20]
  reg  confReg_406; // @[ScanConf.scala 32:20]
  reg  confReg_407; // @[ScanConf.scala 32:20]
  reg  confReg_408; // @[ScanConf.scala 32:20]
  reg  confReg_409; // @[ScanConf.scala 32:20]
  reg  confReg_410; // @[ScanConf.scala 32:20]
  reg  confReg_411; // @[ScanConf.scala 32:20]
  reg  confReg_412; // @[ScanConf.scala 32:20]
  reg  confReg_413; // @[ScanConf.scala 32:20]
  reg  confReg_414; // @[ScanConf.scala 32:20]
  reg  confReg_415; // @[ScanConf.scala 32:20]
  reg  confReg_416; // @[ScanConf.scala 32:20]
  reg  confReg_417; // @[ScanConf.scala 32:20]
  reg  confReg_418; // @[ScanConf.scala 32:20]
  reg  confReg_419; // @[ScanConf.scala 32:20]
  reg  confReg_420; // @[ScanConf.scala 32:20]
  reg  confReg_421; // @[ScanConf.scala 32:20]
  reg  confReg_422; // @[ScanConf.scala 32:20]
  reg  confReg_423; // @[ScanConf.scala 32:20]
  wire [3:0] io_scan_out_lo = {confReg_3,confReg_2,confReg_1,confReg_0}; // @[ScanConf.scala 46:47]
  wire [3:0] io_scan_out_hi = {confReg_7,confReg_6,confReg_5,confReg_4}; // @[ScanConf.scala 46:47]
  wire [5:0] io_confOut_lo_lo_lo_lo_lo_lo = {confReg_5,confReg_4,confReg_3,confReg_2,confReg_1,confReg_0}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_lo_lo_lo_lo_lo = {confReg_12,confReg_11,confReg_10,confReg_9,confReg_8,confReg_7,confReg_6,
    io_confOut_lo_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_lo_lo_lo_hi_lo = {confReg_18,confReg_17,confReg_16,confReg_15,confReg_14,confReg_13}; // @[ScanConf.scala 48:25]
  wire [25:0] io_confOut_lo_lo_lo_lo = {confReg_25,confReg_24,confReg_23,confReg_22,confReg_21,confReg_20,confReg_19,
    io_confOut_lo_lo_lo_lo_hi_lo,io_confOut_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_lo_lo_hi_lo_lo = {confReg_31,confReg_30,confReg_29,confReg_28,confReg_27,confReg_26}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_lo_lo_lo_hi_lo = {confReg_38,confReg_37,confReg_36,confReg_35,confReg_34,confReg_33,confReg_32,
    io_confOut_lo_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_lo_lo_hi_hi_lo = {confReg_45,confReg_44,confReg_43,confReg_42,confReg_41,confReg_40,
    confReg_39}; // @[ScanConf.scala 48:25]
  wire [52:0] io_confOut_lo_lo_lo = {confReg_52,confReg_51,confReg_50,confReg_49,confReg_48,confReg_47,confReg_46,
    io_confOut_lo_lo_lo_hi_hi_lo,io_confOut_lo_lo_lo_hi_lo,io_confOut_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_lo_hi_lo_lo_lo = {confReg_58,confReg_57,confReg_56,confReg_55,confReg_54,confReg_53}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_lo_lo_hi_lo_lo = {confReg_65,confReg_64,confReg_63,confReg_62,confReg_61,confReg_60,confReg_59,
    io_confOut_lo_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_lo_hi_lo_hi_lo = {confReg_71,confReg_70,confReg_69,confReg_68,confReg_67,confReg_66}; // @[ScanConf.scala 48:25]
  wire [25:0] io_confOut_lo_lo_hi_lo = {confReg_78,confReg_77,confReg_76,confReg_75,confReg_74,confReg_73,confReg_72,
    io_confOut_lo_lo_hi_lo_hi_lo,io_confOut_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_lo_hi_hi_lo_lo = {confReg_84,confReg_83,confReg_82,confReg_81,confReg_80,confReg_79}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_lo_lo_hi_hi_lo = {confReg_91,confReg_90,confReg_89,confReg_88,confReg_87,confReg_86,confReg_85,
    io_confOut_lo_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_lo_hi_hi_hi_lo = {confReg_98,confReg_97,confReg_96,confReg_95,confReg_94,confReg_93,
    confReg_92}; // @[ScanConf.scala 48:25]
  wire [52:0] io_confOut_lo_lo_hi = {confReg_105,confReg_104,confReg_103,confReg_102,confReg_101,confReg_100,confReg_99,
    io_confOut_lo_lo_hi_hi_hi_lo,io_confOut_lo_lo_hi_hi_lo,io_confOut_lo_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_hi_lo_lo_lo_lo = {confReg_111,confReg_110,confReg_109,confReg_108,confReg_107,confReg_106}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_lo_hi_lo_lo_lo = {confReg_118,confReg_117,confReg_116,confReg_115,confReg_114,confReg_113,
    confReg_112,io_confOut_lo_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_hi_lo_lo_hi_lo = {confReg_124,confReg_123,confReg_122,confReg_121,confReg_120,confReg_119}; // @[ScanConf.scala 48:25]
  wire [25:0] io_confOut_lo_hi_lo_lo = {confReg_131,confReg_130,confReg_129,confReg_128,confReg_127,confReg_126,
    confReg_125,io_confOut_lo_hi_lo_lo_hi_lo,io_confOut_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_hi_lo_hi_lo_lo = {confReg_137,confReg_136,confReg_135,confReg_134,confReg_133,confReg_132}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_lo_hi_lo_hi_lo = {confReg_144,confReg_143,confReg_142,confReg_141,confReg_140,confReg_139,
    confReg_138,io_confOut_lo_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_hi_lo_hi_hi_lo = {confReg_151,confReg_150,confReg_149,confReg_148,confReg_147,confReg_146,
    confReg_145}; // @[ScanConf.scala 48:25]
  wire [52:0] io_confOut_lo_hi_lo = {confReg_158,confReg_157,confReg_156,confReg_155,confReg_154,confReg_153,confReg_152
    ,io_confOut_lo_hi_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi_lo,io_confOut_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_hi_hi_lo_lo_lo = {confReg_164,confReg_163,confReg_162,confReg_161,confReg_160,confReg_159}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_lo_hi_hi_lo_lo = {confReg_171,confReg_170,confReg_169,confReg_168,confReg_167,confReg_166,
    confReg_165,io_confOut_lo_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_hi_hi_lo_hi_lo = {confReg_177,confReg_176,confReg_175,confReg_174,confReg_173,confReg_172}; // @[ScanConf.scala 48:25]
  wire [25:0] io_confOut_lo_hi_hi_lo = {confReg_184,confReg_183,confReg_182,confReg_181,confReg_180,confReg_179,
    confReg_178,io_confOut_lo_hi_hi_lo_hi_lo,io_confOut_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_lo_hi_hi_hi_lo_lo = {confReg_190,confReg_189,confReg_188,confReg_187,confReg_186,confReg_185}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_lo_hi_hi_hi_lo = {confReg_197,confReg_196,confReg_195,confReg_194,confReg_193,confReg_192,
    confReg_191,io_confOut_lo_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_hi_hi_hi_hi_lo = {confReg_204,confReg_203,confReg_202,confReg_201,confReg_200,confReg_199,
    confReg_198}; // @[ScanConf.scala 48:25]
  wire [52:0] io_confOut_lo_hi_hi = {confReg_211,confReg_210,confReg_209,confReg_208,confReg_207,confReg_206,confReg_205
    ,io_confOut_lo_hi_hi_hi_hi_lo,io_confOut_lo_hi_hi_hi_lo,io_confOut_lo_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [211:0] io_confOut_lo = {io_confOut_lo_hi_hi,io_confOut_lo_hi_lo,io_confOut_lo_lo_hi,io_confOut_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_lo_lo_lo_lo_lo = {confReg_217,confReg_216,confReg_215,confReg_214,confReg_213,confReg_212}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_hi_lo_lo_lo_lo = {confReg_224,confReg_223,confReg_222,confReg_221,confReg_220,confReg_219,
    confReg_218,io_confOut_hi_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_lo_lo_lo_hi_lo = {confReg_230,confReg_229,confReg_228,confReg_227,confReg_226,confReg_225}; // @[ScanConf.scala 48:25]
  wire [25:0] io_confOut_hi_lo_lo_lo = {confReg_237,confReg_236,confReg_235,confReg_234,confReg_233,confReg_232,
    confReg_231,io_confOut_hi_lo_lo_lo_hi_lo,io_confOut_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_lo_lo_hi_lo_lo = {confReg_243,confReg_242,confReg_241,confReg_240,confReg_239,confReg_238}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_hi_lo_lo_hi_lo = {confReg_250,confReg_249,confReg_248,confReg_247,confReg_246,confReg_245,
    confReg_244,io_confOut_hi_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_lo_lo_hi_hi_lo = {confReg_257,confReg_256,confReg_255,confReg_254,confReg_253,confReg_252,
    confReg_251}; // @[ScanConf.scala 48:25]
  wire [52:0] io_confOut_hi_lo_lo = {confReg_264,confReg_263,confReg_262,confReg_261,confReg_260,confReg_259,confReg_258
    ,io_confOut_hi_lo_lo_hi_hi_lo,io_confOut_hi_lo_lo_hi_lo,io_confOut_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_lo_hi_lo_lo_lo = {confReg_270,confReg_269,confReg_268,confReg_267,confReg_266,confReg_265}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_hi_lo_hi_lo_lo = {confReg_277,confReg_276,confReg_275,confReg_274,confReg_273,confReg_272,
    confReg_271,io_confOut_hi_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_lo_hi_lo_hi_lo = {confReg_283,confReg_282,confReg_281,confReg_280,confReg_279,confReg_278}; // @[ScanConf.scala 48:25]
  wire [25:0] io_confOut_hi_lo_hi_lo = {confReg_290,confReg_289,confReg_288,confReg_287,confReg_286,confReg_285,
    confReg_284,io_confOut_hi_lo_hi_lo_hi_lo,io_confOut_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_lo_hi_hi_lo_lo = {confReg_296,confReg_295,confReg_294,confReg_293,confReg_292,confReg_291}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_hi_lo_hi_hi_lo = {confReg_303,confReg_302,confReg_301,confReg_300,confReg_299,confReg_298,
    confReg_297,io_confOut_hi_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_lo_hi_hi_hi_lo = {confReg_310,confReg_309,confReg_308,confReg_307,confReg_306,confReg_305,
    confReg_304}; // @[ScanConf.scala 48:25]
  wire [52:0] io_confOut_hi_lo_hi = {confReg_317,confReg_316,confReg_315,confReg_314,confReg_313,confReg_312,confReg_311
    ,io_confOut_hi_lo_hi_hi_hi_lo,io_confOut_hi_lo_hi_hi_lo,io_confOut_hi_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_hi_lo_lo_lo_lo = {confReg_323,confReg_322,confReg_321,confReg_320,confReg_319,confReg_318}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_hi_hi_lo_lo_lo = {confReg_330,confReg_329,confReg_328,confReg_327,confReg_326,confReg_325,
    confReg_324,io_confOut_hi_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_hi_lo_lo_hi_lo = {confReg_336,confReg_335,confReg_334,confReg_333,confReg_332,confReg_331}; // @[ScanConf.scala 48:25]
  wire [25:0] io_confOut_hi_hi_lo_lo = {confReg_343,confReg_342,confReg_341,confReg_340,confReg_339,confReg_338,
    confReg_337,io_confOut_hi_hi_lo_lo_hi_lo,io_confOut_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_hi_lo_hi_lo_lo = {confReg_349,confReg_348,confReg_347,confReg_346,confReg_345,confReg_344}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_hi_hi_lo_hi_lo = {confReg_356,confReg_355,confReg_354,confReg_353,confReg_352,confReg_351,
    confReg_350,io_confOut_hi_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_hi_lo_hi_hi_lo = {confReg_363,confReg_362,confReg_361,confReg_360,confReg_359,confReg_358,
    confReg_357}; // @[ScanConf.scala 48:25]
  wire [52:0] io_confOut_hi_hi_lo = {confReg_370,confReg_369,confReg_368,confReg_367,confReg_366,confReg_365,confReg_364
    ,io_confOut_hi_hi_lo_hi_hi_lo,io_confOut_hi_hi_lo_hi_lo,io_confOut_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_hi_hi_lo_lo_lo = {confReg_376,confReg_375,confReg_374,confReg_373,confReg_372,confReg_371}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_hi_hi_hi_lo_lo = {confReg_383,confReg_382,confReg_381,confReg_380,confReg_379,confReg_378,
    confReg_377,io_confOut_hi_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_hi_hi_lo_hi_lo = {confReg_389,confReg_388,confReg_387,confReg_386,confReg_385,confReg_384}; // @[ScanConf.scala 48:25]
  wire [25:0] io_confOut_hi_hi_hi_lo = {confReg_396,confReg_395,confReg_394,confReg_393,confReg_392,confReg_391,
    confReg_390,io_confOut_hi_hi_hi_lo_hi_lo,io_confOut_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [5:0] io_confOut_hi_hi_hi_hi_lo_lo = {confReg_402,confReg_401,confReg_400,confReg_399,confReg_398,confReg_397}; // @[ScanConf.scala 48:25]
  wire [12:0] io_confOut_hi_hi_hi_hi_lo = {confReg_409,confReg_408,confReg_407,confReg_406,confReg_405,confReg_404,
    confReg_403,io_confOut_hi_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_hi_hi_hi_hi_lo = {confReg_416,confReg_415,confReg_414,confReg_413,confReg_412,confReg_411,
    confReg_410}; // @[ScanConf.scala 48:25]
  wire [52:0] io_confOut_hi_hi_hi = {confReg_423,confReg_422,confReg_421,confReg_420,confReg_419,confReg_418,confReg_417
    ,io_confOut_hi_hi_hi_hi_hi_lo,io_confOut_hi_hi_hi_hi_lo,io_confOut_hi_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [211:0] io_confOut_hi = {io_confOut_hi_hi_hi,io_confOut_hi_hi_lo,io_confOut_hi_lo_hi,io_confOut_hi_lo_lo}; // @[ScanConf.scala 48:25]
  assign ioBundle_confOut = {io_confOut_hi,io_confOut_lo}; // @[ScanConf.scala 48:25]
  assign ioBundle_scan_out = {io_scan_out_hi,io_scan_out_lo}; // @[ScanConf.scala 46:47]
  always @(posedge clock) begin
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_0 <= confReg_8; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_1 <= confReg_9; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_2 <= confReg_10; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_3 <= confReg_11; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_4 <= confReg_12; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_5 <= confReg_13; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_6 <= confReg_14; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_7 <= confReg_15; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_8 <= confReg_16; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_9 <= confReg_17; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_10 <= confReg_18; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_11 <= confReg_19; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_12 <= confReg_20; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_13 <= confReg_21; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_14 <= confReg_22; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_15 <= confReg_23; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_16 <= confReg_24; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_17 <= confReg_25; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_18 <= confReg_26; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_19 <= confReg_27; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_20 <= confReg_28; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_21 <= confReg_29; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_22 <= confReg_30; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_23 <= confReg_31; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_24 <= confReg_32; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_25 <= confReg_33; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_26 <= confReg_34; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_27 <= confReg_35; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_28 <= confReg_36; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_29 <= confReg_37; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_30 <= confReg_38; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_31 <= confReg_39; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_32 <= confReg_40; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_33 <= confReg_41; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_34 <= confReg_42; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_35 <= confReg_43; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_36 <= confReg_44; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_37 <= confReg_45; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_38 <= confReg_46; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_39 <= confReg_47; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_40 <= confReg_48; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_41 <= confReg_49; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_42 <= confReg_50; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_43 <= confReg_51; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_44 <= confReg_52; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_45 <= confReg_53; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_46 <= confReg_54; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_47 <= confReg_55; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_48 <= confReg_56; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_49 <= confReg_57; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_50 <= confReg_58; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_51 <= confReg_59; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_52 <= confReg_60; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_53 <= confReg_61; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_54 <= confReg_62; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_55 <= confReg_63; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_56 <= confReg_64; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_57 <= confReg_65; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_58 <= confReg_66; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_59 <= confReg_67; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_60 <= confReg_68; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_61 <= confReg_69; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_62 <= confReg_70; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_63 <= confReg_71; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_64 <= confReg_72; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_65 <= confReg_73; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_66 <= confReg_74; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_67 <= confReg_75; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_68 <= confReg_76; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_69 <= confReg_77; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_70 <= confReg_78; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_71 <= confReg_79; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_72 <= confReg_80; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_73 <= confReg_81; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_74 <= confReg_82; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_75 <= confReg_83; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_76 <= confReg_84; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_77 <= confReg_85; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_78 <= confReg_86; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_79 <= confReg_87; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_80 <= confReg_88; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_81 <= confReg_89; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_82 <= confReg_90; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_83 <= confReg_91; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_84 <= confReg_92; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_85 <= confReg_93; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_86 <= confReg_94; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_87 <= confReg_95; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_88 <= confReg_96; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_89 <= confReg_97; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_90 <= confReg_98; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_91 <= confReg_99; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_92 <= confReg_100; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_93 <= confReg_101; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_94 <= confReg_102; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_95 <= confReg_103; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_96 <= confReg_104; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_97 <= confReg_105; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_98 <= confReg_106; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_99 <= confReg_107; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_100 <= confReg_108; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_101 <= confReg_109; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_102 <= confReg_110; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_103 <= confReg_111; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_104 <= confReg_112; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_105 <= confReg_113; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_106 <= confReg_114; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_107 <= confReg_115; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_108 <= confReg_116; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_109 <= confReg_117; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_110 <= confReg_118; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_111 <= confReg_119; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_112 <= confReg_120; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_113 <= confReg_121; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_114 <= confReg_122; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_115 <= confReg_123; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_116 <= confReg_124; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_117 <= confReg_125; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_118 <= confReg_126; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_119 <= confReg_127; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_120 <= confReg_128; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_121 <= confReg_129; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_122 <= confReg_130; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_123 <= confReg_131; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_124 <= confReg_132; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_125 <= confReg_133; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_126 <= confReg_134; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_127 <= confReg_135; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_128 <= confReg_136; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_129 <= confReg_137; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_130 <= confReg_138; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_131 <= confReg_139; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_132 <= confReg_140; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_133 <= confReg_141; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_134 <= confReg_142; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_135 <= confReg_143; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_136 <= confReg_144; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_137 <= confReg_145; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_138 <= confReg_146; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_139 <= confReg_147; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_140 <= confReg_148; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_141 <= confReg_149; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_142 <= confReg_150; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_143 <= confReg_151; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_144 <= confReg_152; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_145 <= confReg_153; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_146 <= confReg_154; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_147 <= confReg_155; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_148 <= confReg_156; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_149 <= confReg_157; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_150 <= confReg_158; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_151 <= confReg_159; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_152 <= confReg_160; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_153 <= confReg_161; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_154 <= confReg_162; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_155 <= confReg_163; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_156 <= confReg_164; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_157 <= confReg_165; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_158 <= confReg_166; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_159 <= confReg_167; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_160 <= confReg_168; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_161 <= confReg_169; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_162 <= confReg_170; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_163 <= confReg_171; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_164 <= confReg_172; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_165 <= confReg_173; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_166 <= confReg_174; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_167 <= confReg_175; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_168 <= confReg_176; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_169 <= confReg_177; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_170 <= confReg_178; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_171 <= confReg_179; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_172 <= confReg_180; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_173 <= confReg_181; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_174 <= confReg_182; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_175 <= confReg_183; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_176 <= confReg_184; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_177 <= confReg_185; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_178 <= confReg_186; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_179 <= confReg_187; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_180 <= confReg_188; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_181 <= confReg_189; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_182 <= confReg_190; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_183 <= confReg_191; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_184 <= confReg_192; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_185 <= confReg_193; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_186 <= confReg_194; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_187 <= confReg_195; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_188 <= confReg_196; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_189 <= confReg_197; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_190 <= confReg_198; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_191 <= confReg_199; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_192 <= confReg_200; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_193 <= confReg_201; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_194 <= confReg_202; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_195 <= confReg_203; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_196 <= confReg_204; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_197 <= confReg_205; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_198 <= confReg_206; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_199 <= confReg_207; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_200 <= confReg_208; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_201 <= confReg_209; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_202 <= confReg_210; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_203 <= confReg_211; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_204 <= confReg_212; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_205 <= confReg_213; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_206 <= confReg_214; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_207 <= confReg_215; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_208 <= confReg_216; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_209 <= confReg_217; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_210 <= confReg_218; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_211 <= confReg_219; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_212 <= confReg_220; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_213 <= confReg_221; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_214 <= confReg_222; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_215 <= confReg_223; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_216 <= confReg_224; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_217 <= confReg_225; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_218 <= confReg_226; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_219 <= confReg_227; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_220 <= confReg_228; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_221 <= confReg_229; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_222 <= confReg_230; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_223 <= confReg_231; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_224 <= confReg_232; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_225 <= confReg_233; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_226 <= confReg_234; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_227 <= confReg_235; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_228 <= confReg_236; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_229 <= confReg_237; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_230 <= confReg_238; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_231 <= confReg_239; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_232 <= confReg_240; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_233 <= confReg_241; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_234 <= confReg_242; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_235 <= confReg_243; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_236 <= confReg_244; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_237 <= confReg_245; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_238 <= confReg_246; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_239 <= confReg_247; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_240 <= confReg_248; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_241 <= confReg_249; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_242 <= confReg_250; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_243 <= confReg_251; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_244 <= confReg_252; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_245 <= confReg_253; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_246 <= confReg_254; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_247 <= confReg_255; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_248 <= confReg_256; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_249 <= confReg_257; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_250 <= confReg_258; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_251 <= confReg_259; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_252 <= confReg_260; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_253 <= confReg_261; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_254 <= confReg_262; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_255 <= confReg_263; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_256 <= confReg_264; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_257 <= confReg_265; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_258 <= confReg_266; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_259 <= confReg_267; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_260 <= confReg_268; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_261 <= confReg_269; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_262 <= confReg_270; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_263 <= confReg_271; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_264 <= confReg_272; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_265 <= confReg_273; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_266 <= confReg_274; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_267 <= confReg_275; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_268 <= confReg_276; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_269 <= confReg_277; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_270 <= confReg_278; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_271 <= confReg_279; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_272 <= confReg_280; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_273 <= confReg_281; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_274 <= confReg_282; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_275 <= confReg_283; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_276 <= confReg_284; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_277 <= confReg_285; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_278 <= confReg_286; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_279 <= confReg_287; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_280 <= confReg_288; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_281 <= confReg_289; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_282 <= confReg_290; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_283 <= confReg_291; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_284 <= confReg_292; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_285 <= confReg_293; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_286 <= confReg_294; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_287 <= confReg_295; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_288 <= confReg_296; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_289 <= confReg_297; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_290 <= confReg_298; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_291 <= confReg_299; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_292 <= confReg_300; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_293 <= confReg_301; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_294 <= confReg_302; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_295 <= confReg_303; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_296 <= confReg_304; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_297 <= confReg_305; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_298 <= confReg_306; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_299 <= confReg_307; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_300 <= confReg_308; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_301 <= confReg_309; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_302 <= confReg_310; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_303 <= confReg_311; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_304 <= confReg_312; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_305 <= confReg_313; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_306 <= confReg_314; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_307 <= confReg_315; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_308 <= confReg_316; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_309 <= confReg_317; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_310 <= confReg_318; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_311 <= confReg_319; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_312 <= confReg_320; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_313 <= confReg_321; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_314 <= confReg_322; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_315 <= confReg_323; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_316 <= confReg_324; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_317 <= confReg_325; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_318 <= confReg_326; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_319 <= confReg_327; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_320 <= confReg_328; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_321 <= confReg_329; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_322 <= confReg_330; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_323 <= confReg_331; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_324 <= confReg_332; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_325 <= confReg_333; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_326 <= confReg_334; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_327 <= confReg_335; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_328 <= confReg_336; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_329 <= confReg_337; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_330 <= confReg_338; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_331 <= confReg_339; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_332 <= confReg_340; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_333 <= confReg_341; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_334 <= confReg_342; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_335 <= confReg_343; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_336 <= confReg_344; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_337 <= confReg_345; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_338 <= confReg_346; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_339 <= confReg_347; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_340 <= confReg_348; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_341 <= confReg_349; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_342 <= confReg_350; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_343 <= confReg_351; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_344 <= confReg_352; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_345 <= confReg_353; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_346 <= confReg_354; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_347 <= confReg_355; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_348 <= confReg_356; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_349 <= confReg_357; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_350 <= confReg_358; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_351 <= confReg_359; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_352 <= confReg_360; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_353 <= confReg_361; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_354 <= confReg_362; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_355 <= confReg_363; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_356 <= confReg_364; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_357 <= confReg_365; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_358 <= confReg_366; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_359 <= confReg_367; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_360 <= confReg_368; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_361 <= confReg_369; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_362 <= confReg_370; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_363 <= confReg_371; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_364 <= confReg_372; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_365 <= confReg_373; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_366 <= confReg_374; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_367 <= confReg_375; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_368 <= confReg_376; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_369 <= confReg_377; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_370 <= confReg_378; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_371 <= confReg_379; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_372 <= confReg_380; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_373 <= confReg_381; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_374 <= confReg_382; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_375 <= confReg_383; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_376 <= confReg_384; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_377 <= confReg_385; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_378 <= confReg_386; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_379 <= confReg_387; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_380 <= confReg_388; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_381 <= confReg_389; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_382 <= confReg_390; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_383 <= confReg_391; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_384 <= confReg_392; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_385 <= confReg_393; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_386 <= confReg_394; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_387 <= confReg_395; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_388 <= confReg_396; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_389 <= confReg_397; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_390 <= confReg_398; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_391 <= confReg_399; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_392 <= confReg_400; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_393 <= confReg_401; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_394 <= confReg_402; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_395 <= confReg_403; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_396 <= confReg_404; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_397 <= confReg_405; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_398 <= confReg_406; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_399 <= confReg_407; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_400 <= confReg_408; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_401 <= confReg_409; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_402 <= confReg_410; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_403 <= confReg_411; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_404 <= confReg_412; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_405 <= confReg_413; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_406 <= confReg_414; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_407 <= confReg_415; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_408 <= confReg_416; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_409 <= confReg_417; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_410 <= confReg_418; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_411 <= confReg_419; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_412 <= confReg_420; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_413 <= confReg_421; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_414 <= confReg_422; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_415 <= confReg_423; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_416 <= ioBundle_scan_in[0]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_417 <= ioBundle_scan_in[1]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_418 <= ioBundle_scan_in[2]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_419 <= ioBundle_scan_in[3]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_420 <= ioBundle_scan_in[4]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_421 <= ioBundle_scan_in[5]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_422 <= ioBundle_scan_in[6]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_423 <= ioBundle_scan_in[7]; // @[ScanConf.scala 38:72]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  confReg_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  confReg_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  confReg_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  confReg_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  confReg_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  confReg_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  confReg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  confReg_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  confReg_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  confReg_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  confReg_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  confReg_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  confReg_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  confReg_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  confReg_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  confReg_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  confReg_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  confReg_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  confReg_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  confReg_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  confReg_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  confReg_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  confReg_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  confReg_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  confReg_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  confReg_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  confReg_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  confReg_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  confReg_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  confReg_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  confReg_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  confReg_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  confReg_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  confReg_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  confReg_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  confReg_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  confReg_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  confReg_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  confReg_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  confReg_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  confReg_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  confReg_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  confReg_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  confReg_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  confReg_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  confReg_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  confReg_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  confReg_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  confReg_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  confReg_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  confReg_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  confReg_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  confReg_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  confReg_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  confReg_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  confReg_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  confReg_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  confReg_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  confReg_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  confReg_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  confReg_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  confReg_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  confReg_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  confReg_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  confReg_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  confReg_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  confReg_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  confReg_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  confReg_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  confReg_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  confReg_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  confReg_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  confReg_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  confReg_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  confReg_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  confReg_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  confReg_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  confReg_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  confReg_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  confReg_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  confReg_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  confReg_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  confReg_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  confReg_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  confReg_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  confReg_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  confReg_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  confReg_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  confReg_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  confReg_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  confReg_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  confReg_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  confReg_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  confReg_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  confReg_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  confReg_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  confReg_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  confReg_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  confReg_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  confReg_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  confReg_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  confReg_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  confReg_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  confReg_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  confReg_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  confReg_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  confReg_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  confReg_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  confReg_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  confReg_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  confReg_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  confReg_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  confReg_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  confReg_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  confReg_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  confReg_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  confReg_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  confReg_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  confReg_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  confReg_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  confReg_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  confReg_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  confReg_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  confReg_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  confReg_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  confReg_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  confReg_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  confReg_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  confReg_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  confReg_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  confReg_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  confReg_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  confReg_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  confReg_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  confReg_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  confReg_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  confReg_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  confReg_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  confReg_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  confReg_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  confReg_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  confReg_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  confReg_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  confReg_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  confReg_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  confReg_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  confReg_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  confReg_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  confReg_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  confReg_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  confReg_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  confReg_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  confReg_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  confReg_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  confReg_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  confReg_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  confReg_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  confReg_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  confReg_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  confReg_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  confReg_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  confReg_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  confReg_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  confReg_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  confReg_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  confReg_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  confReg_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  confReg_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  confReg_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  confReg_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  confReg_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  confReg_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  confReg_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  confReg_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  confReg_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  confReg_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  confReg_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  confReg_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  confReg_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  confReg_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  confReg_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  confReg_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  confReg_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  confReg_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  confReg_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  confReg_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  confReg_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  confReg_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  confReg_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  confReg_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  confReg_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  confReg_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  confReg_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  confReg_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  confReg_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  confReg_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  confReg_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  confReg_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  confReg_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  confReg_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  confReg_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  confReg_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  confReg_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  confReg_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  confReg_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  confReg_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  confReg_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  confReg_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  confReg_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  confReg_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  confReg_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  confReg_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  confReg_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  confReg_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  confReg_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  confReg_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  confReg_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  confReg_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  confReg_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  confReg_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  confReg_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  confReg_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  confReg_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  confReg_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  confReg_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  confReg_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  confReg_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  confReg_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  confReg_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  confReg_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  confReg_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  confReg_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  confReg_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  confReg_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  confReg_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  confReg_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  confReg_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  confReg_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  confReg_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  confReg_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  confReg_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  confReg_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  confReg_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  confReg_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  confReg_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  confReg_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  confReg_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  confReg_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  confReg_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  confReg_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  confReg_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  confReg_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  confReg_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  confReg_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  confReg_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  confReg_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  confReg_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  confReg_257 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  confReg_258 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  confReg_259 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  confReg_260 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  confReg_261 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  confReg_262 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  confReg_263 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  confReg_264 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  confReg_265 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  confReg_266 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  confReg_267 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  confReg_268 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  confReg_269 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  confReg_270 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  confReg_271 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  confReg_272 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  confReg_273 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  confReg_274 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  confReg_275 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  confReg_276 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  confReg_277 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  confReg_278 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  confReg_279 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  confReg_280 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  confReg_281 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  confReg_282 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  confReg_283 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  confReg_284 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  confReg_285 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  confReg_286 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  confReg_287 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  confReg_288 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  confReg_289 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  confReg_290 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  confReg_291 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  confReg_292 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  confReg_293 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  confReg_294 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  confReg_295 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  confReg_296 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  confReg_297 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  confReg_298 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  confReg_299 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  confReg_300 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  confReg_301 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  confReg_302 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  confReg_303 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  confReg_304 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  confReg_305 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  confReg_306 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  confReg_307 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  confReg_308 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  confReg_309 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  confReg_310 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  confReg_311 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  confReg_312 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  confReg_313 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  confReg_314 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  confReg_315 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  confReg_316 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  confReg_317 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  confReg_318 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  confReg_319 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  confReg_320 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  confReg_321 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  confReg_322 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  confReg_323 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  confReg_324 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  confReg_325 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  confReg_326 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  confReg_327 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  confReg_328 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  confReg_329 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  confReg_330 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  confReg_331 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  confReg_332 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  confReg_333 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  confReg_334 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  confReg_335 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  confReg_336 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  confReg_337 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  confReg_338 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  confReg_339 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  confReg_340 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  confReg_341 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  confReg_342 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  confReg_343 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  confReg_344 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  confReg_345 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  confReg_346 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  confReg_347 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  confReg_348 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  confReg_349 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  confReg_350 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  confReg_351 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  confReg_352 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  confReg_353 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  confReg_354 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  confReg_355 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  confReg_356 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  confReg_357 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  confReg_358 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  confReg_359 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  confReg_360 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  confReg_361 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  confReg_362 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  confReg_363 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  confReg_364 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  confReg_365 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  confReg_366 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  confReg_367 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  confReg_368 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  confReg_369 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  confReg_370 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  confReg_371 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  confReg_372 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  confReg_373 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  confReg_374 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  confReg_375 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  confReg_376 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  confReg_377 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  confReg_378 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  confReg_379 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  confReg_380 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  confReg_381 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  confReg_382 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  confReg_383 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  confReg_384 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  confReg_385 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  confReg_386 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  confReg_387 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  confReg_388 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  confReg_389 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  confReg_390 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  confReg_391 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  confReg_392 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  confReg_393 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  confReg_394 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  confReg_395 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  confReg_396 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  confReg_397 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  confReg_398 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  confReg_399 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  confReg_400 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  confReg_401 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  confReg_402 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  confReg_403 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  confReg_404 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  confReg_405 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  confReg_406 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  confReg_407 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  confReg_408 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  confReg_409 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  confReg_410 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  confReg_411 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  confReg_412 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  confReg_413 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  confReg_414 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  confReg_415 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  confReg_416 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  confReg_417 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  confReg_418 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  confReg_419 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  confReg_420 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  confReg_421 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  confReg_422 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  confReg_423 = _RAND_423[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MuxNInput_18_SCAOptCB(
  input  [17:0] io_in,
  input  [4:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [31:0] OPinMux_in; // @[MuxListTest.scala 44:28]
  wire [4:0] OPinMux_sel; // @[MuxListTest.scala 44:28]
  wire  OPinMux_o; // @[MuxListTest.scala 44:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux32C OPinMux ( // @[MuxListTest.scala 44:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{14'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_16_SCAOptCB(
  input  [15:0] io_in,
  input  [4:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [31:0] OPinMux_in; // @[MuxListTest.scala 44:28]
  wire [4:0] OPinMux_sel; // @[MuxListTest.scala 44:28]
  wire  OPinMux_o; // @[MuxListTest.scala 44:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux32C OPinMux ( // @[MuxListTest.scala 44:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{16'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_20_SCAOptCB(
  input  [19:0] io_in,
  input  [4:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [31:0] OPinMux_in; // @[MuxListTest.scala 44:28]
  wire [4:0] OPinMux_sel; // @[MuxListTest.scala 44:28]
  wire  OPinMux_o; // @[MuxListTest.scala 44:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux32C OPinMux ( // @[MuxListTest.scala 44:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{12'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_O7_C1_SCAOptSB(
  input  [7:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{1'd0}, io_in[6:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{7'd0}, io_in[7]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O6_C1_SCAOptSB(
  input  [6:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{2'd0}, io_in[5:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{7'd0}, io_in[6]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O6_C2_SCAOptSB(
  input  [7:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{2'd0}, io_in[5:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{6'd0}, io_in[7:6]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O7_C2_SCAOptSB(
  input  [8:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{1'd0}, io_in[6:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{6'd0}, io_in[8:7]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O16_C1_SCAOptSB(
  input  [16:0] io_in,
  input  [4:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_ioGndBle,
  input         io_cnstClk,
  input         io_arst
);
  wire [15:0] OPinMux_in; // @[MuxListTest.scala 111:26]
  wire [3:0] OPinMux_sel; // @[MuxListTest.scala 111:26]
  wire  OPinMux_o; // @[MuxListTest.scala 111:26]
  wire [15:0] chanMux_in; // @[MuxListTest.scala 132:26]
  wire [3:0] chanMux_sel; // @[MuxListTest.scala 132:26]
  wire  chanMux_o; // @[MuxListTest.scala 132:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux16C OPinMux ( // @[MuxListTest.scala 111:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux16C chanMux ( // @[MuxListTest.scala 132:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = io_in[15:0]; // @[MuxListTest.scala 123:30]
  assign OPinMux_sel = io_config[3:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{15'd0}, io_in[16]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[3:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[4] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O0_C5_SCAOptSB(
  input  [4:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = 8'h0; // @[MuxListTest.scala 125:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module Tile_11_3_iotile(
  input          clock,
  input          reset,
  input          IN_OPIN_N22321_33,
  input          IN_OPIN_N22323_35,
  input          IN_OPIN_N22325_37,
  input          IN_OPIN_N22327_39,
  input          IN_OPIN_N22329_41,
  input          IN_OPIN_N22331_43,
  input          IN_OPIN_N22333_45,
  input          IN_OPIN_N22335_47,
  input          IN_OPIN_N22337_49,
  input          IN_OPIN_N22339_51,
  input          IN_OPIN_N22341_53,
  input          IN_OPIN_N22343_55,
  input          IN_OPIN_N22345_57,
  input          IN_OPIN_N22347_59,
  input          IN_OPIN_N22349_61,
  input          IN_OPIN_N22351_63,
  input          IN_CHANX_N24196_4,
  input          IN_CHANX_N24198_12,
  input          IN_CHANX_N24200_20,
  input          IN_CHANX_N24202_28,
  input          IN_CHANX_N24204_36,
  input          IN_CHANX_N24206_44,
  input          IN_CHANX_N24208_52,
  input          IN_CHANX_N24210_60,
  input          IN_CHANX_N24212_68,
  input          IN_CHANX_N24216_6,
  input          IN_CHANX_N24218_14,
  input          IN_CHANX_N24220_22,
  input          IN_CHANX_N24222_30,
  input          IN_CHANX_N24224_38,
  input          IN_CHANX_N24226_46,
  input          IN_CHANX_N24228_54,
  input          IN_CHANX_N24230_62,
  input          IN_CHANX_N24232_70,
  input          IN_CHANX_N24236_0,
  input          IN_CHANX_N24238_8,
  input          IN_CHANX_N24240_16,
  input          IN_CHANX_N24242_24,
  input          IN_CHANX_N24244_32,
  input          IN_CHANX_N24246_40,
  input          IN_CHANX_N24248_48,
  input          IN_CHANX_N24250_56,
  input          IN_CHANX_N24252_64,
  input          IN_CHANX_N24254_72,
  input          IN_CHANX_N24256_76,
  input          IN_CHANX_N24258_2,
  input          IN_CHANX_N24260_10,
  input          IN_CHANX_N24262_18,
  input          IN_CHANX_N24264_26,
  input          IN_CHANX_N24266_34,
  input          IN_CHANX_N24268_42,
  input          IN_CHANX_N24270_50,
  input          IN_CHANX_N24272_58,
  input          IN_CHANX_N24274_66,
  input          IN_CHANX_N24276_74,
  input          IN_CHANX_N24278_78,
  input          IN_CHANY_N29000_2,
  input          IN_CHANY_N29001_3,
  input          IN_CHANY_N29002_4,
  input          IN_CHANY_N29003_5,
  input          IN_CHANY_N29008_10,
  input          IN_CHANY_N29009_11,
  input          IN_CHANY_N29010_12,
  input          IN_CHANY_N29011_13,
  input          IN_CHANY_N29016_18,
  input          IN_CHANY_N29017_19,
  input          IN_CHANY_N29018_20,
  input          IN_CHANY_N29019_21,
  input          IN_CHANY_N29024_26,
  input          IN_CHANY_N29025_27,
  input          IN_CHANY_N29026_28,
  input          IN_CHANY_N29027_29,
  input          IN_CHANY_N29032_34,
  input          IN_CHANY_N29033_35,
  input          IN_CHANY_N29034_36,
  input          IN_CHANY_N29035_37,
  input          IN_CHANY_N29078_6,
  input          IN_CHANY_N29079_7,
  input          IN_CHANY_N29080_14,
  input          IN_CHANY_N29081_15,
  input          IN_CHANY_N29082_22,
  input          IN_CHANY_N29083_23,
  input          IN_CHANY_N29084_30,
  input          IN_CHANY_N29085_31,
  input          IN_CHANY_N29096_78,
  input          IN_CHANY_N29097_79,
  input          IN_CHANY_N29098_0,
  input          IN_CHANY_N29099_1,
  input          IN_CHANY_N29100_8,
  input          IN_CHANY_N29101_9,
  input          IN_CHANY_N29102_16,
  input          IN_CHANY_N29103_17,
  input          IN_CHANY_N29104_24,
  input          IN_CHANY_N29105_25,
  input          IN_CHANY_N29106_32,
  input          IN_CHANY_N29107_33,
  input          IN_CHANY_N29108_40,
  input          IN_CHANY_N29109_41,
  input          IN_CHANY_N29110_48,
  input          IN_CHANY_N29111_49,
  input          IN_CHANY_N29112_56,
  input          IN_CHANY_N29113_57,
  input          IN_CHANY_N29114_64,
  input          IN_CHANY_N29115_65,
  input          IN_CHANY_N29116_72,
  input          IN_CHANY_N29117_73,
  input          IN_CHANY_N29118_76,
  input          IN_CHANY_N29119_77,
  input          IN_CHANY_N29270_4,
  input          IN_CHANY_N29272_6,
  input          IN_CHANY_N29273_7,
  input          IN_CHANY_N29278_12,
  input          IN_CHANY_N29280_14,
  input          IN_CHANY_N29281_15,
  input          IN_CHANY_N29286_20,
  input          IN_CHANY_N29288_22,
  input          IN_CHANY_N29289_23,
  input          IN_CHANY_N29294_28,
  input          IN_CHANY_N29296_30,
  input          IN_CHANY_N29297_31,
  input          IN_CHANY_N29302_36,
  input          IN_CHANY_N29310_44,
  input          IN_CHANY_N29318_52,
  input          IN_CHANY_N29326_60,
  input          IN_CHANY_N29334_68,
  input          IN_CHANY_N29346_0,
  input          IN_CHANY_N29347_1,
  input          IN_CHANY_N29348_8,
  input          IN_CHANY_N29349_9,
  input          IN_CHANY_N29350_16,
  input          IN_CHANY_N29351_17,
  input          IN_CHANY_N29352_24,
  input          IN_CHANY_N29353_25,
  input          IN_CHANY_N29354_32,
  input          IN_CHANY_N29355_33,
  input          IN_CHANY_N29366_76,
  input          IN_CHANY_N29368_2,
  input          IN_CHANY_N29369_3,
  input          IN_CHANY_N29370_10,
  input          IN_CHANY_N29371_11,
  input          IN_CHANY_N29372_18,
  input          IN_CHANY_N29373_19,
  input          IN_CHANY_N29374_26,
  input          IN_CHANY_N29375_27,
  input          IN_CHANY_N29376_34,
  input          IN_CHANY_N29377_35,
  input          IN_CHANY_N29378_42,
  input          IN_CHANY_N29379_43,
  input          IN_CHANY_N29380_50,
  input          IN_CHANY_N29381_51,
  input          IN_CHANY_N29382_58,
  input          IN_CHANY_N29383_59,
  input          IN_CHANY_N29384_66,
  input          IN_CHANY_N29385_67,
  input          IN_CHANY_N29386_74,
  input          IN_CHANY_N29387_75,
  input          IN_CHANY_N29388_78,
  input          IN_CHANY_N29389_79,
  input          IN_CHANY_N29391_5,
  input          IN_CHANY_N29393_13,
  input          IN_CHANY_N29395_21,
  input          IN_CHANY_N29397_29,
  input          IN_CHANY_N29399_37,
  input          IN_CHANY_N29401_45,
  input          IN_CHANY_N29403_53,
  input          IN_CHANY_N29405_61,
  input          IN_CHANY_N29407_69,
  input          IN_CHANY_N29409_77,
  output         OUT_OPIN_N22211_51,
  output         OUT_CHANY_N29400_44,
  output         OUT_CHANX_N24229_55,
  output         OUT_CHANX_N24239_9,
  output         OUT_CHANX_N24269_43,
  output         OUT_CHANY_N29398_36,
  output         OUT_CHANX_N24237_1,
  output         OUT_CHANX_N24199_13,
  output         OUT_CHANX_N24211_61,
  output         OUT_OPIN_N22223_63,
  output         OUT_CHANX_N24241_17,
  output         OUT_CHANX_N24213_69,
  output         OUT_CHANX_N24279_79,
  output         OUT_OPIN_N22193_33,
  output         OUT_CHANX_N24207_45,
  output         OUT_OPIN_N22185_25,
  output         OUT_CHANX_N24233_71,
  output         OUT_CHANX_N24221_23,
  output         OUT_CHANX_N24271_51,
  output         OUT_OPIN_N22187_27,
  output         OUT_CHANX_N24245_33,
  output         OUT_CHANX_N24265_27,
  output         OUT_CHANY_N29390_4,
  output         OUT_CHANY_N29319_53,
  output         OUT_CHANX_N24209_53,
  output         OUT_CHANX_N24217_7,
  output         OUT_CHANX_N24273_59,
  output         OUT_CHANY_N29408_76,
  output         OUT_CHANY_N29287_21,
  output         OUT_CHANX_N24197_5,
  output         OUT_CHANX_N24267_35,
  output         OUT_CHANX_N24203_29,
  output         OUT_OPIN_N22183_23,
  output         OUT_CHANY_N29271_5,
  output         OUT_CHANY_N29406_68,
  output         OUT_CHANX_N24219_15,
  output         OUT_OPIN_N22161_1,
  output         OUT_CHANX_N24201_21,
  output         OUT_OPIN_N22215_55,
  output         OUT_CHANX_N24253_65,
  output         OUT_CHANY_N29295_29,
  output         OUT_OPIN_N22175_15,
  output         OUT_OPIN_N22217_57,
  output         OUT_OPIN_N22213_53,
  output         OUT_CHANY_N29303_37,
  output         OUT_CHANY_N29311_45,
  output         OUT_OPIN_N22177_17,
  output         OUT_CHANY_N29392_12,
  output         OUT_CHANX_N24205_37,
  output         OUT_CHANX_N24247_41,
  output         OUT_OPIN_N22163_3,
  output         OUT_OPIN_N22165_5,
  output         OUT_OPIN_N22189_29,
  output         OUT_CHANX_N24255_73,
  output         OUT_CHANX_N24263_19,
  output         OUT_OPIN_N22169_9,
  output         OUT_OPIN_N22207_47,
  output         OUT_OPIN_N22201_41,
  output         OUT_OPIN_N22205_45,
  output         OUT_CHANX_N24251_57,
  output         OUT_OPIN_N22219_59,
  output         OUT_CHANY_N29402_52,
  output         OUT_CHANY_N29367_77,
  output         OUT_CHANY_N29394_20,
  output         OUT_CHANX_N24259_3,
  output         OUT_OPIN_N22221_61,
  output         OUT_CHANX_N24223_31,
  output         OUT_CHANX_N24231_63,
  output         OUT_OPIN_N22181_21,
  output         OUT_CHANY_N29404_60,
  output         OUT_CHANY_N29327_61,
  output         OUT_OPIN_N22171_11,
  output         OUT_CHANX_N24261_11,
  output         OUT_OPIN_N22195_35,
  output         OUT_OPIN_N22179_19,
  output         OUT_CHANX_N24275_67,
  output         OUT_CHANY_N29396_28,
  output         OUT_CHANX_N24243_25,
  output         OUT_OPIN_N22167_7,
  output         OUT_OPIN_N22197_37,
  output         OUT_OPIN_N22209_49,
  output         OUT_CHANY_N29279_13,
  output         OUT_CHANX_N24277_75,
  output         OUT_OPIN_N22199_39,
  output         OUT_CHANX_N24249_49,
  output         OUT_OPIN_N22203_43,
  output         OUT_OPIN_N22173_13,
  output         OUT_CHANY_N29335_69,
  output         OUT_CHANX_N24227_47,
  output         OUT_CHANX_N24257_77,
  output         OUT_CHANX_N24225_39,
  output         OUT_OPIN_N22191_31,
  output [417:0] ioConf_confOut,
  input  [7:0]   ioConf_scan_in,
  input          ioConf_scan_en,
  output [7:0]   ioConf_scan_out,
  input  [31:0]  ioPad_i,
  output [31:0]  ioPad_o,
  input          ctrlSignals_gndBlkOuts,
  input          ctrlSignals_loopBreak,
  input          ctrlSignals_arst,
  input          ctrlSignals_tmrMode,
  input          ctrlSignals_confClock,
  input          ctrlSignals_constClock
);
  wire  logicBlock_IPIN_0; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_2; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_4; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_6; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_8; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_10; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_12; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_14; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_16; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_18; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_20; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_22; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_24; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_26; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_28; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_30; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_32; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_34; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_36; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_38; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_40; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_42; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_44; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_46; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_48; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_50; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_52; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_54; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_56; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_58; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_60; // @[TileFull.scala 44:33]
  wire  logicBlock_IPIN_62; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_1; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_3; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_5; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_7; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_9; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_11; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_13; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_15; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_17; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_19; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_21; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_23; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_25; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_27; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_29; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_31; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_33; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_35; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_37; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_39; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_41; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_43; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_45; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_47; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_49; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_51; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_53; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_55; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_57; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_59; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_61; // @[TileFull.scala 44:33]
  wire  logicBlock_OPIN_63; // @[TileFull.scala 44:33]
  wire  logicBlock_clock; // @[TileFull.scala 44:33]
  wire  logicBlock_reset; // @[TileFull.scala 44:33]
  wire [31:0] logicBlock_ioPad_i; // @[TileFull.scala 44:33]
  wire [31:0] logicBlock_ioPad_o; // @[TileFull.scala 44:33]
  wire [15:0] logicBlock_configBits; // @[TileFull.scala 44:33]
  wire  logicBlock_loopBreak; // @[TileFull.scala 44:33]
  wire  logicBlock_gndLBouts; // @[TileFull.scala 44:33]
  wire  configBlock_clock; // @[TileFull.scala 61:31]
  wire [423:0] configBlock_ioBundle_confOut; // @[TileFull.scala 61:31]
  wire [7:0] configBlock_ioBundle_scan_in; // @[TileFull.scala 61:31]
  wire  configBlock_ioBundle_scan_en; // @[TileFull.scala 61:31]
  wire [7:0] configBlock_ioBundle_scan_out; // @[TileFull.scala 61:31]
  wire [17:0] CBMux_IPIN0_N22160_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN0_N22160_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N22160_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N22160_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N22160_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N22160_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN2_N22162_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN2_N22162_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N22162_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N22162_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N22162_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N22162_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN4_N22164_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN4_N22164_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N22164_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N22164_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N22164_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N22164_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN6_N22166_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN6_N22166_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N22166_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N22166_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N22166_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N22166_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN8_N22168_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN8_N22168_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N22168_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N22168_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N22168_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N22168_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN10_N22170_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN10_N22170_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N22170_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N22170_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N22170_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N22170_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN12_N22172_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN12_N22172_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N22172_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N22172_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N22172_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N22172_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN14_N22174_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN14_N22174_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N22174_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N22174_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N22174_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N22174_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN16_N22176_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN16_N22176_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N22176_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N22176_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N22176_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N22176_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN18_N22178_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN18_N22178_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N22178_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N22178_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N22178_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N22178_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN20_N22180_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN20_N22180_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N22180_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N22180_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N22180_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N22180_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN22_N22182_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN22_N22182_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N22182_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N22182_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N22182_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N22182_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN24_N22184_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN24_N22184_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N22184_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N22184_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N22184_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N22184_io_arst; // @[TileFull.scala 97:27]
  wire [19:0] CBMux_IPIN26_N22186_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN26_N22186_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N22186_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N22186_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N22186_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N22186_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN28_N22188_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN28_N22188_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N22188_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N22188_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N22188_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N22188_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN30_N22190_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN30_N22190_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N22190_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N22190_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N22190_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N22190_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN32_N22192_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN32_N22192_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N22192_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N22192_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N22192_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N22192_io_arst; // @[TileFull.scala 97:27]
  wire [19:0] CBMux_IPIN34_N22194_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN34_N22194_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N22194_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N22194_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N22194_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N22194_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN36_N22196_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN36_N22196_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N22196_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N22196_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N22196_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N22196_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN38_N22198_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN38_N22198_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N22198_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N22198_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N22198_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N22198_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN40_N22200_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN40_N22200_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN40_N22200_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN40_N22200_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN40_N22200_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN40_N22200_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN42_N22202_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN42_N22202_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN42_N22202_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN42_N22202_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN42_N22202_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN42_N22202_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN44_N22204_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN44_N22204_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN44_N22204_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN44_N22204_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN44_N22204_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN44_N22204_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN46_N22206_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN46_N22206_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN46_N22206_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN46_N22206_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN46_N22206_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN46_N22206_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN48_N22208_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN48_N22208_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN48_N22208_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN48_N22208_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN48_N22208_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN48_N22208_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN50_N22210_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN50_N22210_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN50_N22210_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN50_N22210_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN50_N22210_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN50_N22210_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN52_N22212_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN52_N22212_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN52_N22212_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN52_N22212_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN52_N22212_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN52_N22212_io_arst; // @[TileFull.scala 97:27]
  wire [15:0] CBMux_IPIN54_N22214_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN54_N22214_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN54_N22214_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN54_N22214_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN54_N22214_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN54_N22214_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN56_N22216_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN56_N22216_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN56_N22216_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN56_N22216_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN56_N22216_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN56_N22216_io_arst; // @[TileFull.scala 97:27]
  wire [19:0] CBMux_IPIN58_N22218_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN58_N22218_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN58_N22218_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN58_N22218_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN58_N22218_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN58_N22218_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN60_N22220_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN60_N22220_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN60_N22220_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN60_N22220_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN60_N22220_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN60_N22220_io_arst; // @[TileFull.scala 97:27]
  wire [17:0] CBMux_IPIN62_N22222_io_in; // @[TileFull.scala 97:27]
  wire [4:0] CBMux_IPIN62_N22222_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN62_N22222_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN62_N22222_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN62_N22222_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN62_N22222_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] SBMux_C5_N24197_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C5_N24197_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N24197_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N24197_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N24197_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N24197_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N24197_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C13_N24199_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C13_N24199_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N24199_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N24199_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N24199_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N24199_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N24199_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C21_N24201_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C21_N24201_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N24201_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N24201_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N24201_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N24201_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N24201_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [6:0] SBMux_C29_N24203_O_6_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C29_N24203_O_6_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N24203_O_6_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N24203_O_6_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N24203_O_6_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N24203_O_6_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N24203_O_6_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C37_N24205_O_6_C_2_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C37_N24205_O_6_C_2_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N24205_O_6_C_2_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N24205_O_6_C_2_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N24205_O_6_C_2_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N24205_O_6_C_2_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N24205_O_6_C_2_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C45_N24207_O_7_C_2_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C45_N24207_O_7_C_2_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N24207_O_7_C_2_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N24207_O_7_C_2_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N24207_O_7_C_2_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N24207_O_7_C_2_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N24207_O_7_C_2_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C53_N24209_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C53_N24209_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N24209_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N24209_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N24209_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N24209_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N24209_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C61_N24211_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C61_N24211_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N24211_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N24211_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N24211_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N24211_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N24211_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [6:0] SBMux_C69_N24213_O_6_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C69_N24213_O_6_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N24213_O_6_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N24213_O_6_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N24213_O_6_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N24213_O_6_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N24213_O_6_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C7_N24217_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C7_N24217_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C7_N24217_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C7_N24217_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C7_N24217_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C7_N24217_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C7_N24217_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C15_N24219_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C15_N24219_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C15_N24219_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C15_N24219_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C15_N24219_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C15_N24219_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C15_N24219_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C23_N24221_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C23_N24221_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C23_N24221_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C23_N24221_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C23_N24221_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C23_N24221_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C23_N24221_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [6:0] SBMux_C31_N24223_O_6_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C31_N24223_O_6_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C31_N24223_O_6_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C31_N24223_O_6_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C31_N24223_O_6_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C31_N24223_O_6_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C31_N24223_O_6_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C39_N24225_O_7_C_2_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C39_N24225_O_7_C_2_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C39_N24225_O_7_C_2_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C39_N24225_O_7_C_2_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C39_N24225_O_7_C_2_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C39_N24225_O_7_C_2_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C39_N24225_O_7_C_2_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C47_N24227_O_7_C_2_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C47_N24227_O_7_C_2_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C47_N24227_O_7_C_2_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C47_N24227_O_7_C_2_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C47_N24227_O_7_C_2_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C47_N24227_O_7_C_2_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C47_N24227_O_7_C_2_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C55_N24229_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C55_N24229_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C55_N24229_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C55_N24229_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C55_N24229_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C55_N24229_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C55_N24229_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C63_N24231_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C63_N24231_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C63_N24231_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C63_N24231_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C63_N24231_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C63_N24231_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C63_N24231_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [6:0] SBMux_C71_N24233_O_6_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C71_N24233_O_6_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C71_N24233_O_6_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C71_N24233_O_6_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C71_N24233_O_6_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C71_N24233_O_6_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C71_N24233_O_6_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C1_N24237_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C1_N24237_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N24237_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N24237_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N24237_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N24237_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N24237_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C9_N24239_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C9_N24239_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N24239_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N24239_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N24239_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N24239_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N24239_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C17_N24241_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C17_N24241_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N24241_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N24241_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N24241_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N24241_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N24241_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C25_N24243_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C25_N24243_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N24243_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N24243_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N24243_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N24243_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N24243_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [6:0] SBMux_C33_N24245_O_6_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C33_N24245_O_6_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N24245_O_6_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N24245_O_6_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N24245_O_6_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N24245_O_6_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N24245_O_6_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C41_N24247_O_7_C_2_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C41_N24247_O_7_C_2_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N24247_O_7_C_2_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N24247_O_7_C_2_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N24247_O_7_C_2_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N24247_O_7_C_2_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N24247_O_7_C_2_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C49_N24249_O_7_C_2_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C49_N24249_O_7_C_2_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N24249_O_7_C_2_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N24249_O_7_C_2_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N24249_O_7_C_2_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N24249_O_7_C_2_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N24249_O_7_C_2_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C57_N24251_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C57_N24251_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N24251_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N24251_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N24251_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N24251_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N24251_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C65_N24253_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C65_N24253_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N24253_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N24253_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N24253_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N24253_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N24253_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [6:0] SBMux_C73_N24255_O_6_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C73_N24255_O_6_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N24255_O_6_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N24255_O_6_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N24255_O_6_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N24255_O_6_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N24255_O_6_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [16:0] SBMux_C77_N24257_O_16_C_1_io_in; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C77_N24257_O_16_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24257_O_16_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24257_O_16_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24257_O_16_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24257_O_16_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24257_O_16_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C3_N24259_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C3_N24259_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C3_N24259_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C3_N24259_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C3_N24259_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C3_N24259_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C3_N24259_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C11_N24261_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C11_N24261_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C11_N24261_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C11_N24261_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C11_N24261_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C11_N24261_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C11_N24261_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C19_N24263_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C19_N24263_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C19_N24263_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C19_N24263_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C19_N24263_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C19_N24263_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C19_N24263_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C27_N24265_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C27_N24265_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C27_N24265_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C27_N24265_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C27_N24265_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C27_N24265_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C27_N24265_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C35_N24267_O_6_C_2_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C35_N24267_O_6_C_2_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C35_N24267_O_6_C_2_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C35_N24267_O_6_C_2_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C35_N24267_O_6_C_2_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C35_N24267_O_6_C_2_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C35_N24267_O_6_C_2_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C43_N24269_O_7_C_2_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C43_N24269_O_7_C_2_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C43_N24269_O_7_C_2_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C43_N24269_O_7_C_2_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C43_N24269_O_7_C_2_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C43_N24269_O_7_C_2_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C43_N24269_O_7_C_2_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C51_N24271_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C51_N24271_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C51_N24271_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C51_N24271_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C51_N24271_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C51_N24271_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C51_N24271_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C59_N24273_O_7_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C59_N24273_O_7_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C59_N24273_O_7_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C59_N24273_O_7_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C59_N24273_O_7_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C59_N24273_O_7_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C59_N24273_O_7_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [6:0] SBMux_C67_N24275_O_6_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C67_N24275_O_6_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C67_N24275_O_6_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C67_N24275_O_6_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C67_N24275_O_6_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C67_N24275_O_6_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C67_N24275_O_6_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [6:0] SBMux_C75_N24277_O_6_C_1_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C75_N24277_O_6_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C75_N24277_O_6_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C75_N24277_O_6_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C75_N24277_O_6_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C75_N24277_O_6_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C75_N24277_O_6_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [16:0] SBMux_C79_N24279_O_16_C_1_io_in; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C79_N24279_O_16_C_1_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C79_N24279_O_16_C_1_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C79_N24279_O_16_C_1_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C79_N24279_O_16_C_1_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C79_N24279_O_16_C_1_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C79_N24279_O_16_C_1_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C5_N29271_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C5_N29271_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N29271_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N29271_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N29271_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N29271_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C5_N29271_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C13_N29279_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C13_N29279_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N29279_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N29279_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N29279_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N29279_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C13_N29279_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C21_N29287_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C21_N29287_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N29287_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N29287_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N29287_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N29287_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C21_N29287_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C29_N29295_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C29_N29295_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N29295_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N29295_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N29295_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N29295_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C29_N29295_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C37_N29303_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C37_N29303_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N29303_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N29303_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N29303_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N29303_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C37_N29303_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C45_N29311_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C45_N29311_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N29311_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N29311_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N29311_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N29311_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C45_N29311_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C53_N29319_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C53_N29319_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N29319_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N29319_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N29319_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N29319_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C53_N29319_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C61_N29327_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C61_N29327_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N29327_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N29327_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N29327_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N29327_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C61_N29327_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C69_N29335_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C69_N29335_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N29335_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N29335_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N29335_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N29335_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C69_N29335_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C77_N29367_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C77_N29367_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N29367_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N29367_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N29367_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N29367_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N29367_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C4_N29390_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C4_N29390_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N29390_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N29390_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N29390_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N29390_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C4_N29390_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C12_N29392_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C12_N29392_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N29392_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N29392_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N29392_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N29392_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C12_N29392_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C20_N29394_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C20_N29394_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N29394_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N29394_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N29394_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N29394_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C20_N29394_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C28_N29396_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C28_N29396_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N29396_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N29396_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N29396_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N29396_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C28_N29396_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C36_N29398_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C36_N29398_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N29398_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N29398_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N29398_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N29398_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C36_N29398_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C44_N29400_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C44_N29400_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N29400_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N29400_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N29400_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N29400_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C44_N29400_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C52_N29402_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C52_N29402_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N29402_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N29402_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N29402_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N29402_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C52_N29402_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C60_N29404_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C60_N29404_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N29404_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N29404_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N29404_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N29404_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C60_N29404_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C68_N29406_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C68_N29406_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N29406_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N29406_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N29406_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N29406_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C68_N29406_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] SBMux_C76_N29408_O_0_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C76_N29408_O_0_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N29408_O_0_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N29408_O_0_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N29408_O_0_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N29408_O_0_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N29408_O_0_C_5_io_arst; // @[TileFull.scala 134:27]
  wire  _CBMux_IPIN0_N22160_io_in_WIRE_1 = SBMux_C5_N29271_O_0_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN0_N22160_io_in_WIRE_5 = SBMux_C29_N29295_O_0_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [8:0] CBMux_IPIN0_N22160_io_in_lo = {IN_CHANY_N29350_16,IN_CHANY_N29297_31,IN_CHANY_N29296_30,
    _CBMux_IPIN0_N22160_io_in_WIRE_5,IN_CHANY_N29294_28,IN_CHANY_N29273_7,IN_CHANY_N29272_6,
    _CBMux_IPIN0_N22160_io_in_WIRE_1,IN_CHANY_N29270_4}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN0_N22160_io_in_hi = {IN_CHANY_N29389_79,IN_CHANY_N29388_78,IN_CHANY_N29385_67,IN_CHANY_N29384_66,
    IN_CHANY_N29379_43,IN_CHANY_N29378_42,IN_CHANY_N29371_11,IN_CHANY_N29370_10,IN_CHANY_N29351_17}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN2_N22162_io_in_WIRE_1 = SBMux_C13_N29279_O_0_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN2_N22162_io_in_WIRE_5 = SBMux_C37_N29303_O_0_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [8:0] CBMux_IPIN2_N22162_io_in_lo = {IN_CHANY_N29352_24,IN_CHANY_N29347_1,IN_CHANY_N29346_0,
    _CBMux_IPIN2_N22162_io_in_WIRE_5,IN_CHANY_N29302_36,IN_CHANY_N29281_15,IN_CHANY_N29280_14,
    _CBMux_IPIN2_N22162_io_in_WIRE_1,IN_CHANY_N29278_12}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN2_N22162_io_in_WIRE_11 = SBMux_C77_N29367_O_0_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [8:0] CBMux_IPIN2_N22162_io_in_hi = {IN_CHANY_N29387_75,IN_CHANY_N29386_74,IN_CHANY_N29381_51,IN_CHANY_N29380_50,
    IN_CHANY_N29373_19,IN_CHANY_N29372_18,_CBMux_IPIN2_N22162_io_in_WIRE_11,IN_CHANY_N29366_76,IN_CHANY_N29353_25}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN4_N22164_io_in_WIRE_1 = SBMux_C21_N29287_O_0_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [7:0] CBMux_IPIN4_N22164_io_in_lo = {IN_CHANY_N29355_33,IN_CHANY_N29354_32,IN_CHANY_N29349_9,IN_CHANY_N29348_8,
    IN_CHANY_N29289_23,IN_CHANY_N29288_22,_CBMux_IPIN4_N22164_io_in_WIRE_1,IN_CHANY_N29286_20}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN4_N22164_io_in_hi = {IN_CHANY_N29383_59,IN_CHANY_N29382_58,IN_CHANY_N29375_27,IN_CHANY_N29374_26,
    IN_CHANY_N29369_3,IN_CHANY_N29368_2,_CBMux_IPIN2_N22162_io_in_WIRE_11,IN_CHANY_N29366_76}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN6_N22166_io_in_lo = {IN_CHANY_N29369_3,IN_CHANY_N29368_2,IN_CHANY_N29349_9,IN_CHANY_N29348_8,
    IN_CHANY_N29289_23,IN_CHANY_N29288_22,_CBMux_IPIN4_N22164_io_in_WIRE_1,IN_CHANY_N29286_20}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN6_N22166_io_in_hi = {IN_CHANY_N29389_79,IN_CHANY_N29388_78,IN_CHANY_N29383_59,IN_CHANY_N29382_58,
    IN_CHANY_N29377_35,IN_CHANY_N29376_34,IN_CHANY_N29375_27,IN_CHANY_N29374_26}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN8_N22168_io_in_lo = {IN_CHANY_N29350_16,_CBMux_IPIN2_N22162_io_in_WIRE_5,IN_CHANY_N29302_36,
    IN_CHANY_N29297_31,IN_CHANY_N29296_30,IN_CHANY_N29273_7,IN_CHANY_N29272_6,_CBMux_IPIN0_N22160_io_in_WIRE_1,
    IN_CHANY_N29270_4}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN8_N22168_io_in_hi = {IN_CHANY_N29389_79,IN_CHANY_N29388_78,IN_CHANY_N29387_75,IN_CHANY_N29386_74,
    IN_CHANY_N29379_43,IN_CHANY_N29378_42,IN_CHANY_N29371_11,IN_CHANY_N29370_10,IN_CHANY_N29351_17}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN10_N22170_io_in_lo = {IN_CHANY_N29353_25,IN_CHANY_N29352_24,IN_CHANY_N29347_1,IN_CHANY_N29346_0,
    IN_CHANY_N29281_15,IN_CHANY_N29280_14,_CBMux_IPIN2_N22162_io_in_WIRE_1,IN_CHANY_N29278_12}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN10_N22170_io_in_hi = {IN_CHANY_N29381_51,IN_CHANY_N29380_50,IN_CHANY_N29373_19,IN_CHANY_N29372_18
    ,_CBMux_IPIN2_N22162_io_in_WIRE_11,IN_CHANY_N29366_76,IN_CHANY_N29355_33,IN_CHANY_N29354_32}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN12_N22172_io_in_lo = {IN_CHANY_N29366_76,IN_CHANY_N29349_9,IN_CHANY_N29348_8,
    _CBMux_IPIN0_N22160_io_in_WIRE_5,IN_CHANY_N29294_28,IN_CHANY_N29289_23,IN_CHANY_N29288_22,
    _CBMux_IPIN4_N22164_io_in_WIRE_1,IN_CHANY_N29286_20}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN12_N22172_io_in_hi = {IN_CHANY_N29385_67,IN_CHANY_N29384_66,IN_CHANY_N29383_59,IN_CHANY_N29382_58
    ,IN_CHANY_N29377_35,IN_CHANY_N29376_34,IN_CHANY_N29369_3,IN_CHANY_N29368_2,_CBMux_IPIN2_N22162_io_in_WIRE_11}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN14_N22174_io_in_lo = {IN_CHANY_N29370_10,IN_CHANY_N29351_17,IN_CHANY_N29350_16,IN_CHANY_N29297_31
    ,IN_CHANY_N29296_30,_CBMux_IPIN0_N22160_io_in_WIRE_5,IN_CHANY_N29294_28,_CBMux_IPIN0_N22160_io_in_WIRE_1,
    IN_CHANY_N29270_4}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN14_N22174_io_in_hi = {IN_CHANY_N29389_79,IN_CHANY_N29388_78,IN_CHANY_N29385_67,IN_CHANY_N29384_66
    ,IN_CHANY_N29379_43,IN_CHANY_N29378_42,IN_CHANY_N29377_35,IN_CHANY_N29376_34,IN_CHANY_N29371_11}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN16_N22176_io_in_lo = {IN_CHANY_N29352_24,_CBMux_IPIN2_N22162_io_in_WIRE_5,IN_CHANY_N29302_36,
    IN_CHANY_N29281_15,IN_CHANY_N29280_14,_CBMux_IPIN2_N22162_io_in_WIRE_1,IN_CHANY_N29278_12,IN_CHANY_N29273_7,
    IN_CHANY_N29272_6}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN16_N22176_io_in_hi = {IN_CHANY_N29389_79,IN_CHANY_N29388_78,IN_CHANY_N29387_75,IN_CHANY_N29386_74
    ,IN_CHANY_N29381_51,IN_CHANY_N29380_50,IN_CHANY_N29373_19,IN_CHANY_N29372_18,IN_CHANY_N29353_25}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN18_N22178_io_in_lo = {IN_CHANY_N29355_33,IN_CHANY_N29354_32,IN_CHANY_N29347_1,IN_CHANY_N29346_0,
    IN_CHANY_N29281_15,IN_CHANY_N29280_14,_CBMux_IPIN2_N22162_io_in_WIRE_1,IN_CHANY_N29278_12}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN18_N22178_io_in_hi = {IN_CHANY_N29381_51,IN_CHANY_N29380_50,IN_CHANY_N29375_27,IN_CHANY_N29374_26
    ,IN_CHANY_N29373_19,IN_CHANY_N29372_18,_CBMux_IPIN2_N22162_io_in_WIRE_11,IN_CHANY_N29366_76}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN20_N22180_io_in_lo = {IN_CHANY_N29349_9,IN_CHANY_N29348_8,IN_CHANY_N29347_1,IN_CHANY_N29346_0,
    IN_CHANY_N29289_23,IN_CHANY_N29288_22,_CBMux_IPIN4_N22164_io_in_WIRE_1,IN_CHANY_N29286_20}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN20_N22180_io_in_hi = {IN_CHANY_N29383_59,IN_CHANY_N29382_58,IN_CHANY_N29375_27,IN_CHANY_N29374_26
    ,_CBMux_IPIN2_N22162_io_in_WIRE_11,IN_CHANY_N29366_76,IN_CHANY_N29355_33,IN_CHANY_N29354_32}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN22_N22182_io_in_lo = {IN_CHANY_N29369_3,IN_CHANY_N29368_2,IN_CHANY_N29351_17,IN_CHANY_N29350_16,
    IN_CHANY_N29297_31,IN_CHANY_N29296_30,_CBMux_IPIN0_N22160_io_in_WIRE_5,IN_CHANY_N29294_28}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN22_N22182_io_in_hi = {IN_CHANY_N29389_79,IN_CHANY_N29388_78,IN_CHANY_N29385_67,IN_CHANY_N29384_66
    ,IN_CHANY_N29377_35,IN_CHANY_N29376_34,IN_CHANY_N29371_11,IN_CHANY_N29370_10}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN24_N22184_io_in_lo = {IN_CHANY_N29352_24,IN_CHANY_N29351_17,IN_CHANY_N29350_16,
    _CBMux_IPIN2_N22162_io_in_WIRE_5,IN_CHANY_N29302_36,IN_CHANY_N29273_7,IN_CHANY_N29272_6,
    _CBMux_IPIN0_N22160_io_in_WIRE_1,IN_CHANY_N29270_4}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN24_N22184_io_in_hi = {IN_CHANY_N29389_79,IN_CHANY_N29388_78,IN_CHANY_N29387_75,IN_CHANY_N29386_74
    ,IN_CHANY_N29379_43,IN_CHANY_N29378_42,IN_CHANY_N29371_11,IN_CHANY_N29370_10,IN_CHANY_N29353_25}; // @[TileFull.scala 166:8]
  wire [9:0] CBMux_IPIN26_N22186_io_in_lo = {IN_CHANY_N29353_25,IN_CHANY_N29352_24,_CBMux_IPIN2_N22162_io_in_WIRE_5,
    IN_CHANY_N29302_36,_CBMux_IPIN2_N22162_io_in_WIRE_1,IN_CHANY_N29278_12,IN_CHANY_N29273_7,IN_CHANY_N29272_6,
    _CBMux_IPIN0_N22160_io_in_WIRE_1,IN_CHANY_N29270_4}; // @[TileFull.scala 166:8]
  wire [9:0] CBMux_IPIN26_N22186_io_in_hi = {IN_CHANY_N29387_75,IN_CHANY_N29386_74,IN_CHANY_N29381_51,IN_CHANY_N29380_50
    ,IN_CHANY_N29379_43,IN_CHANY_N29378_42,IN_CHANY_N29373_19,IN_CHANY_N29372_18,_CBMux_IPIN2_N22162_io_in_WIRE_11,
    IN_CHANY_N29366_76}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN28_N22188_io_in_lo = {IN_CHANY_N29347_1,IN_CHANY_N29346_0,IN_CHANY_N29289_23,IN_CHANY_N29288_22,
    _CBMux_IPIN4_N22164_io_in_WIRE_1,IN_CHANY_N29286_20,IN_CHANY_N29281_15,IN_CHANY_N29280_14}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN30_N22190_io_in_lo = {IN_CHANY_N29349_9,IN_CHANY_N29348_8,IN_CHANY_N29297_31,IN_CHANY_N29296_30,
    _CBMux_IPIN0_N22160_io_in_WIRE_5,IN_CHANY_N29294_28,IN_CHANY_N29289_23,IN_CHANY_N29288_22}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN30_N22190_io_in_hi = {IN_CHANY_N29389_79,IN_CHANY_N29388_78,IN_CHANY_N29385_67,IN_CHANY_N29384_66
    ,IN_CHANY_N29377_35,IN_CHANY_N29376_34,IN_CHANY_N29369_3,IN_CHANY_N29368_2}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN32_N22192_io_in_lo = {IN_CHANY_N29085_31,IN_CHANY_N29084_30,IN_CHANY_N29079_7,IN_CHANY_N29078_6,
    IN_CHANY_N29017_19,IN_CHANY_N29016_18,IN_CHANY_N29011_13,IN_CHANY_N29010_12}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN32_N22192_io_in_hi = {IN_CHANY_N29119_77,IN_CHANY_N29118_76,IN_CHANY_N29113_57,IN_CHANY_N29112_56
    ,IN_CHANY_N29105_25,IN_CHANY_N29104_24,IN_CHANY_N29099_1,IN_CHANY_N29098_0}; // @[TileFull.scala 166:8]
  wire [9:0] CBMux_IPIN34_N22194_io_in_lo = {IN_CHANY_N29081_15,IN_CHANY_N29080_14,IN_CHANY_N29033_35,IN_CHANY_N29032_34
    ,IN_CHANY_N29025_27,IN_CHANY_N29024_26,IN_CHANY_N29019_21,IN_CHANY_N29018_20,IN_CHANY_N29001_3,IN_CHANY_N29000_2}; // @[TileFull.scala 166:8]
  wire [9:0] CBMux_IPIN34_N22194_io_in_hi = {IN_CHANY_N29117_73,IN_CHANY_N29116_72,IN_CHANY_N29115_65,IN_CHANY_N29114_64
    ,IN_CHANY_N29109_41,IN_CHANY_N29108_40,IN_CHANY_N29101_9,IN_CHANY_N29100_8,IN_CHANY_N29097_79,IN_CHANY_N29096_78}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN36_N22196_io_in_lo = {IN_CHANY_N29035_37,IN_CHANY_N29034_36,IN_CHANY_N29027_29,IN_CHANY_N29026_28
    ,IN_CHANY_N29009_11,IN_CHANY_N29008_10,IN_CHANY_N29003_5,IN_CHANY_N29002_4}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN36_N22196_io_in_hi = {IN_CHANY_N29111_49,IN_CHANY_N29110_48,IN_CHANY_N29103_17,IN_CHANY_N29102_16
    ,IN_CHANY_N29097_79,IN_CHANY_N29096_78,IN_CHANY_N29083_23,IN_CHANY_N29082_22}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN38_N22198_io_in_lo = {IN_CHANY_N29099_1,IN_CHANY_N29098_0,IN_CHANY_N29079_7,IN_CHANY_N29078_6,
    IN_CHANY_N29017_19,IN_CHANY_N29016_18,IN_CHANY_N29011_13,IN_CHANY_N29010_12}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN38_N22198_io_in_hi = {IN_CHANY_N29119_77,IN_CHANY_N29118_76,IN_CHANY_N29113_57,IN_CHANY_N29112_56
    ,IN_CHANY_N29107_33,IN_CHANY_N29106_32,IN_CHANY_N29105_25,IN_CHANY_N29104_24}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN40_N22200_io_in_lo = {IN_CHANY_N29100_8,IN_CHANY_N29081_15,IN_CHANY_N29080_14,IN_CHANY_N29025_27,
    IN_CHANY_N29024_26,IN_CHANY_N29019_21,IN_CHANY_N29018_20,IN_CHANY_N29001_3,IN_CHANY_N29000_2}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN40_N22200_io_in_hi = {IN_CHANY_N29119_77,IN_CHANY_N29118_76,IN_CHANY_N29115_65,IN_CHANY_N29114_64
    ,IN_CHANY_N29109_41,IN_CHANY_N29108_40,IN_CHANY_N29107_33,IN_CHANY_N29106_32,IN_CHANY_N29101_9}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN42_N22202_io_in_lo = {IN_CHANY_N29082_22,IN_CHANY_N29033_35,IN_CHANY_N29032_34,IN_CHANY_N29027_29
    ,IN_CHANY_N29026_28,IN_CHANY_N29009_11,IN_CHANY_N29008_10,IN_CHANY_N29003_5,IN_CHANY_N29002_4}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN42_N22202_io_in_hi = {IN_CHANY_N29117_73,IN_CHANY_N29116_72,IN_CHANY_N29111_49,IN_CHANY_N29110_48
    ,IN_CHANY_N29103_17,IN_CHANY_N29102_16,IN_CHANY_N29097_79,IN_CHANY_N29096_78,IN_CHANY_N29083_23}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN44_N22204_io_in_lo = {IN_CHANY_N29083_23,IN_CHANY_N29082_22,IN_CHANY_N29035_37,IN_CHANY_N29034_36
    ,IN_CHANY_N29009_11,IN_CHANY_N29008_10,IN_CHANY_N29003_5,IN_CHANY_N29002_4}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN44_N22204_io_in_hi = {IN_CHANY_N29111_49,IN_CHANY_N29110_48,IN_CHANY_N29103_17,IN_CHANY_N29102_16
    ,IN_CHANY_N29097_79,IN_CHANY_N29096_78,IN_CHANY_N29085_31,IN_CHANY_N29084_30}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN50_N22210_io_in_lo = {IN_CHANY_N29080_14,IN_CHANY_N29033_35,IN_CHANY_N29032_34,IN_CHANY_N29027_29
    ,IN_CHANY_N29026_28,IN_CHANY_N29019_21,IN_CHANY_N29018_20,IN_CHANY_N29001_3,IN_CHANY_N29000_2}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN50_N22210_io_in_hi = {IN_CHANY_N29117_73,IN_CHANY_N29116_72,IN_CHANY_N29109_41,IN_CHANY_N29108_40
    ,IN_CHANY_N29101_9,IN_CHANY_N29100_8,IN_CHANY_N29097_79,IN_CHANY_N29096_78,IN_CHANY_N29081_15}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN54_N22214_io_in_lo = {IN_CHANY_N29079_7,IN_CHANY_N29078_6,IN_CHANY_N29035_37,IN_CHANY_N29034_36,
    IN_CHANY_N29017_19,IN_CHANY_N29016_18,IN_CHANY_N29011_13,IN_CHANY_N29010_12}; // @[TileFull.scala 166:8]
  wire [7:0] CBMux_IPIN54_N22214_io_in_hi = {IN_CHANY_N29119_77,IN_CHANY_N29118_76,IN_CHANY_N29113_57,IN_CHANY_N29112_56
    ,IN_CHANY_N29105_25,IN_CHANY_N29104_24,IN_CHANY_N29085_31,IN_CHANY_N29084_30}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN56_N22216_io_in_lo = {IN_CHANY_N29098_0,IN_CHANY_N29079_7,IN_CHANY_N29078_6,IN_CHANY_N29025_27,
    IN_CHANY_N29024_26,IN_CHANY_N29017_19,IN_CHANY_N29016_18,IN_CHANY_N29011_13,IN_CHANY_N29010_12}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN56_N22216_io_in_hi = {IN_CHANY_N29119_77,IN_CHANY_N29118_76,IN_CHANY_N29115_65,IN_CHANY_N29114_64
    ,IN_CHANY_N29113_57,IN_CHANY_N29112_56,IN_CHANY_N29107_33,IN_CHANY_N29106_32,IN_CHANY_N29099_1}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN62_N22222_io_in_lo = {IN_CHANY_N29084_30,IN_CHANY_N29035_37,IN_CHANY_N29034_36,IN_CHANY_N29017_19
    ,IN_CHANY_N29016_18,IN_CHANY_N29009_11,IN_CHANY_N29008_10,IN_CHANY_N29003_5,IN_CHANY_N29002_4}; // @[TileFull.scala 166:8]
  wire [8:0] CBMux_IPIN62_N22222_io_in_hi = {IN_CHANY_N29119_77,IN_CHANY_N29118_76,IN_CHANY_N29113_57,IN_CHANY_N29112_56
    ,IN_CHANY_N29111_49,IN_CHANY_N29110_48,IN_CHANY_N29105_25,IN_CHANY_N29104_24,IN_CHANY_N29085_31}; // @[TileFull.scala 166:8]
  wire  _SBMux_C5_N24197_O_7_C_1_io_in_WIRE_1 = logicBlock_OPIN_11; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C5_N24197_O_7_C_1_io_in_WIRE_0 = logicBlock_OPIN_1; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C5_N24197_O_7_C_1_io_in_WIRE_3 = logicBlock_OPIN_29; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C5_N24197_O_7_C_1_io_in_WIRE_2 = logicBlock_OPIN_21; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C5_N24197_O_7_C_1_io_in_lo = {_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_3,
    _SBMux_C5_N24197_O_7_C_1_io_in_WIRE_2,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_1,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C5_N24197_O_7_C_1_io_in_hi = {IN_CHANY_N29278_12,IN_OPIN_N22347_59,IN_OPIN_N22337_49,
    IN_OPIN_N22327_39}; // @[TileFull.scala 183:11]
  wire  _SBMux_C13_N24199_O_7_C_1_io_in_WIRE_1 = logicBlock_OPIN_13; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C13_N24199_O_7_C_1_io_in_WIRE_0 = logicBlock_OPIN_3; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C13_N24199_O_7_C_1_io_in_WIRE_3 = logicBlock_OPIN_31; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C13_N24199_O_7_C_1_io_in_WIRE_2 = logicBlock_OPIN_23; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C13_N24199_O_7_C_1_io_in_lo = {_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_3,
    _SBMux_C13_N24199_O_7_C_1_io_in_WIRE_2,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_1,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_0
    }; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C13_N24199_O_7_C_1_io_in_hi = {IN_CHANY_N29310_44,IN_OPIN_N22349_61,IN_OPIN_N22339_51,
    IN_OPIN_N22329_41}; // @[TileFull.scala 183:11]
  wire  _SBMux_C21_N24201_O_7_C_1_io_in_WIRE_1 = logicBlock_OPIN_15; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C21_N24201_O_7_C_1_io_in_WIRE_0 = logicBlock_OPIN_5; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C21_N24201_O_7_C_1_io_in_WIRE_2 = logicBlock_OPIN_25; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C21_N24201_O_7_C_1_io_in_lo = {IN_OPIN_N22321_33,_SBMux_C21_N24201_O_7_C_1_io_in_WIRE_2,
    _SBMux_C21_N24201_O_7_C_1_io_in_WIRE_1,_SBMux_C21_N24201_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C21_N24201_O_7_C_1_io_in_hi = {IN_CHANY_N29366_76,IN_OPIN_N22351_63,IN_OPIN_N22341_53,
    IN_OPIN_N22331_43}; // @[TileFull.scala 183:11]
  wire  _SBMux_C29_N24203_O_6_C_1_io_in_WIRE_2 = logicBlock_OPIN_27; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C29_N24203_O_6_C_1_io_in_WIRE_1 = logicBlock_OPIN_17; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C29_N24203_O_6_C_1_io_in_WIRE_0 = logicBlock_OPIN_7; // @[TileFull.scala 174:{37,37}]
  wire [2:0] SBMux_C29_N24203_O_6_C_1_io_in_lo = {_SBMux_C29_N24203_O_6_C_1_io_in_WIRE_2,
    _SBMux_C29_N24203_O_6_C_1_io_in_WIRE_1,_SBMux_C29_N24203_O_6_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C29_N24203_O_6_C_1_io_in_hi = {IN_CHANY_N29348_8,IN_OPIN_N22343_55,IN_OPIN_N22333_45,
    IN_OPIN_N22323_35}; // @[TileFull.scala 183:11]
  wire  _SBMux_C37_N24205_O_6_C_2_io_in_WIRE_1 = logicBlock_OPIN_19; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C37_N24205_O_6_C_2_io_in_WIRE_0 = logicBlock_OPIN_9; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C37_N24205_O_6_C_2_io_in_lo = {IN_OPIN_N22325_37,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_3,
    _SBMux_C37_N24205_O_6_C_2_io_in_WIRE_1,_SBMux_C37_N24205_O_6_C_2_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C37_N24205_O_6_C_2_io_in_hi = {IN_CHANY_N29372_18,IN_CHANY_N29355_33,IN_OPIN_N22345_57,
    IN_OPIN_N22335_47}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C45_N24207_O_7_C_2_io_in_lo = {_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_3,
    _SBMux_C5_N24197_O_7_C_1_io_in_WIRE_2,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_1,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C45_N24207_O_7_C_2_io_in_hi = {IN_CHANY_N29296_30,IN_CHANY_N29289_23,IN_OPIN_N22347_59,
    IN_OPIN_N22337_49,IN_OPIN_N22327_39}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C53_N24209_O_7_C_1_io_in_lo = {IN_OPIN_N22321_33,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_2,
    _SBMux_C13_N24199_O_7_C_1_io_in_WIRE_1,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C53_N24209_O_7_C_1_io_in_hi = {IN_CHANY_N29371_11,IN_OPIN_N22349_61,IN_OPIN_N22339_51,
    IN_OPIN_N22329_41}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C61_N24211_O_7_C_1_io_in_lo = {IN_OPIN_N22323_35,_SBMux_C21_N24201_O_7_C_1_io_in_WIRE_2,
    _SBMux_C21_N24201_O_7_C_1_io_in_WIRE_1,_SBMux_C21_N24201_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C61_N24211_O_7_C_1_io_in_hi = {IN_CHANY_N29347_1,IN_OPIN_N22351_63,IN_OPIN_N22341_53,
    IN_OPIN_N22331_43}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C69_N24213_O_6_C_1_io_in_hi = {IN_CHANY_N29403_53,IN_OPIN_N22343_55,IN_OPIN_N22333_45,
    IN_OPIN_N22325_37}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C7_N24217_O_7_C_1_io_in_hi = {IN_CHANY_N29286_20,IN_OPIN_N22347_59,IN_OPIN_N22337_49,
    IN_OPIN_N22327_39}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C15_N24219_O_7_C_1_io_in_hi = {IN_CHANY_N29318_52,IN_OPIN_N22349_61,IN_OPIN_N22339_51,
    IN_OPIN_N22329_41}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C23_N24221_O_7_C_1_io_in_hi = {IN_CHANY_N29346_0,IN_OPIN_N22351_63,IN_OPIN_N22341_53,
    IN_OPIN_N22331_43}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C31_N24223_O_6_C_1_io_in_hi = {IN_CHANY_N29370_10,IN_OPIN_N22343_55,IN_OPIN_N22333_45,
    IN_OPIN_N22325_37}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C39_N24225_O_7_C_2_io_in_lo = {_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_3,
    _SBMux_C37_N24205_O_6_C_2_io_in_WIRE_1,_SBMux_C37_N24205_O_6_C_2_io_in_WIRE_0,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_0}
    ; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C39_N24225_O_7_C_2_io_in_hi = {IN_CHANY_N29297_31,IN_CHANY_N29288_22,IN_OPIN_N22345_57,
    IN_OPIN_N22335_47,IN_OPIN_N22327_39}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C47_N24227_O_7_C_2_io_in_lo = {_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_3,
    _SBMux_C5_N24197_O_7_C_1_io_in_WIRE_2,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_1,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C47_N24227_O_7_C_2_io_in_hi = {IN_CHANY_N29373_19,IN_CHANY_N29354_32,IN_OPIN_N22347_59,
    IN_OPIN_N22337_49,IN_OPIN_N22329_41}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C55_N24229_O_7_C_1_io_in_lo = {IN_OPIN_N22321_33,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_2,
    _SBMux_C13_N24199_O_7_C_1_io_in_WIRE_1,_SBMux_C21_N24201_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C55_N24229_O_7_C_1_io_in_hi = {IN_CHANY_N29349_9,IN_OPIN_N22349_61,IN_OPIN_N22339_51,
    IN_OPIN_N22331_43}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C63_N24231_O_7_C_1_io_in_lo = {IN_OPIN_N22323_35,_SBMux_C21_N24201_O_7_C_1_io_in_WIRE_2,
    _SBMux_C21_N24201_O_7_C_1_io_in_WIRE_1,_SBMux_C29_N24203_O_6_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C63_N24231_O_7_C_1_io_in_hi = {IN_CHANY_N29409_77,IN_OPIN_N22351_63,IN_OPIN_N22341_53,
    IN_OPIN_N22333_45}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C71_N24233_O_6_C_1_io_in_lo = {_SBMux_C29_N24203_O_6_C_1_io_in_WIRE_2,
    _SBMux_C29_N24203_O_6_C_1_io_in_WIRE_1,_SBMux_C37_N24205_O_6_C_2_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C71_N24233_O_6_C_1_io_in_hi = {IN_CHANY_N29401_45,IN_OPIN_N22343_55,IN_OPIN_N22335_47,
    IN_OPIN_N22325_37}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C1_N24237_O_7_C_1_io_in_hi = {IN_CHANY_N29391_5,IN_OPIN_N22345_57,IN_OPIN_N22335_47,IN_OPIN_N22327_39
    }; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C9_N24239_O_7_C_1_io_in_hi = {IN_CHANY_N29294_28,IN_OPIN_N22347_59,IN_OPIN_N22337_49,
    IN_OPIN_N22329_41}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C17_N24241_O_7_C_1_io_in_hi = {IN_CHANY_N29326_60,IN_OPIN_N22349_61,IN_OPIN_N22339_51,
    IN_OPIN_N22331_43}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C25_N24243_O_7_C_1_io_in_hi = {IN_CHANY_N29368_2,IN_OPIN_N22351_63,IN_OPIN_N22341_53,
    IN_OPIN_N22333_45}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C33_N24245_O_6_C_1_io_in_hi = {IN_CHANY_N29280_14,IN_OPIN_N22343_55,IN_OPIN_N22335_47,
    IN_OPIN_N22325_37}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C41_N24247_O_7_C_2_io_in_lo = {_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_3,
    _SBMux_C37_N24205_O_6_C_2_io_in_WIRE_1,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_1,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C41_N24247_O_7_C_2_io_in_hi = {IN_CHANY_N29375_27,IN_CHANY_N29352_24,IN_OPIN_N22345_57,
    IN_OPIN_N22337_49,IN_OPIN_N22327_39}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C49_N24249_O_7_C_2_io_in_lo = {_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_3,
    _SBMux_C5_N24197_O_7_C_1_io_in_WIRE_2,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_1,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_0}
    ; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C49_N24249_O_7_C_2_io_in_hi = {IN_CHANY_N29376_34,IN_CHANY_N29351_17,IN_OPIN_N22347_59,
    IN_OPIN_N22339_51,IN_OPIN_N22329_41}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C57_N24251_O_7_C_1_io_in_lo = {IN_OPIN_N22321_33,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_2,
    _SBMux_C21_N24201_O_7_C_1_io_in_WIRE_1,_SBMux_C21_N24201_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C57_N24251_O_7_C_1_io_in_hi = {IN_CHANY_N29273_7,IN_OPIN_N22349_61,IN_OPIN_N22341_53,
    IN_OPIN_N22331_43}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C65_N24253_O_7_C_1_io_in_lo = {IN_OPIN_N22323_35,_SBMux_C21_N24201_O_7_C_1_io_in_WIRE_2,
    _SBMux_C29_N24203_O_6_C_1_io_in_WIRE_1,_SBMux_C29_N24203_O_6_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C65_N24253_O_7_C_1_io_in_hi = {IN_CHANY_N29407_69,IN_OPIN_N22351_63,IN_OPIN_N22343_55,
    IN_OPIN_N22333_45}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C73_N24255_O_6_C_1_io_in_lo = {_SBMux_C29_N24203_O_6_C_1_io_in_WIRE_2,
    _SBMux_C37_N24205_O_6_C_2_io_in_WIRE_1,_SBMux_C37_N24205_O_6_C_2_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C73_N24255_O_6_C_1_io_in_hi = {IN_CHANY_N29399_37,IN_OPIN_N22345_57,IN_OPIN_N22335_47,
    IN_OPIN_N22325_37}; // @[TileFull.scala 183:11]
  wire [7:0] SBMux_C77_N24257_O_16_C_1_io_in_lo = {_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_3,
    _SBMux_C21_N24201_O_7_C_1_io_in_WIRE_2,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_2,_SBMux_C29_N24203_O_6_C_1_io_in_WIRE_1,
    _SBMux_C13_N24199_O_7_C_1_io_in_WIRE_1,_SBMux_C37_N24205_O_6_C_2_io_in_WIRE_0,_SBMux_C21_N24201_O_7_C_1_io_in_WIRE_0
    ,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [8:0] SBMux_C77_N24257_O_16_C_1_io_in_hi = {IN_CHANY_N29395_21,IN_OPIN_N22349_61,IN_OPIN_N22345_57,
    IN_OPIN_N22341_53,IN_OPIN_N22337_49,IN_OPIN_N22333_45,IN_OPIN_N22329_41,IN_OPIN_N22325_37,IN_OPIN_N22321_33}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C3_N24259_O_7_C_1_io_in_hi = {IN_CHANY_N29270_4,IN_OPIN_N22345_57,IN_OPIN_N22337_49,IN_OPIN_N22327_39
    }; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C11_N24261_O_7_C_1_io_in_hi = {IN_CHANY_N29302_36,IN_OPIN_N22347_59,IN_OPIN_N22339_51,
    IN_OPIN_N22329_41}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C19_N24263_O_7_C_1_io_in_hi = {IN_CHANY_N29334_68,IN_OPIN_N22349_61,IN_OPIN_N22341_53,
    IN_OPIN_N22331_43}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C27_N24265_O_7_C_1_io_in_hi = {IN_CHANY_N29272_6,IN_OPIN_N22351_63,IN_OPIN_N22343_55,
    IN_OPIN_N22333_45}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C35_N24267_O_6_C_2_io_in_lo = {IN_OPIN_N22325_37,_SBMux_C29_N24203_O_6_C_1_io_in_WIRE_2,
    _SBMux_C37_N24205_O_6_C_2_io_in_WIRE_1,_SBMux_C37_N24205_O_6_C_2_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C35_N24267_O_6_C_2_io_in_hi = {IN_CHANY_N29377_35,IN_CHANY_N29350_16,IN_OPIN_N22345_57,
    IN_OPIN_N22335_47}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C43_N24269_O_7_C_2_io_in_hi = {IN_CHANY_N29374_26,IN_CHANY_N29353_25,IN_OPIN_N22347_59,
    IN_OPIN_N22337_49,IN_OPIN_N22327_39}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C51_N24271_O_7_C_1_io_in_hi = {IN_CHANY_N29281_15,IN_OPIN_N22349_61,IN_OPIN_N22339_51,
    IN_OPIN_N22329_41}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C59_N24273_O_7_C_1_io_in_hi = {IN_CHANY_N29369_3,IN_OPIN_N22351_63,IN_OPIN_N22341_53,
    IN_OPIN_N22331_43}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C67_N24275_O_6_C_1_io_in_hi = {IN_CHANY_N29405_61,IN_OPIN_N22343_55,IN_OPIN_N22333_45,
    IN_OPIN_N22323_35}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C75_N24277_O_6_C_1_io_in_lo = {_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_3,
    _SBMux_C37_N24205_O_6_C_2_io_in_WIRE_1,_SBMux_C37_N24205_O_6_C_2_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C75_N24277_O_6_C_1_io_in_hi = {IN_CHANY_N29397_29,IN_OPIN_N22345_57,IN_OPIN_N22335_47,
    IN_OPIN_N22325_37}; // @[TileFull.scala 183:11]
  wire [7:0] SBMux_C79_N24279_O_16_C_1_io_in_lo = {_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_3,
    _SBMux_C29_N24203_O_6_C_1_io_in_WIRE_2,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_2,_SBMux_C37_N24205_O_6_C_2_io_in_WIRE_1
    ,_SBMux_C21_N24201_O_7_C_1_io_in_WIRE_1,_SBMux_C5_N24197_O_7_C_1_io_in_WIRE_1,_SBMux_C29_N24203_O_6_C_1_io_in_WIRE_0
    ,_SBMux_C13_N24199_O_7_C_1_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [8:0] SBMux_C79_N24279_O_16_C_1_io_in_hi = {IN_CHANY_N29393_13,IN_OPIN_N22351_63,IN_OPIN_N22347_59,
    IN_OPIN_N22343_55,IN_OPIN_N22339_51,IN_OPIN_N22335_47,IN_OPIN_N22331_43,IN_OPIN_N22327_39,IN_OPIN_N22323_35}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C5_N29271_O_0_C_5_io_in_lo = {IN_CHANX_N24230_62,IN_CHANX_N24220_22}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C5_N29271_O_0_C_5_io_in_hi = {IN_CHANY_N29391_5,IN_CHANX_N24268_42,IN_CHANX_N24258_2}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C13_N29279_O_0_C_5_io_in_lo = {IN_CHANX_N24206_44,IN_CHANX_N24196_4}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C13_N29279_O_0_C_5_io_in_hi = {IN_CHANY_N29393_13,IN_CHANX_N24252_64,IN_CHANX_N24242_24}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C21_N29287_O_0_C_5_io_in_lo = {IN_CHANX_N24226_46,IN_CHANX_N24216_6}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C21_N29287_O_0_C_5_io_in_hi = {IN_CHANY_N29395_21,IN_CHANX_N24274_66,IN_CHANX_N24264_26}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C29_N29295_O_0_C_5_io_in_lo = {IN_CHANX_N24212_68,IN_CHANX_N24202_28}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C29_N29295_O_0_C_5_io_in_hi = {IN_CHANY_N29397_29,IN_CHANX_N24248_48,IN_CHANX_N24238_8}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C37_N29303_O_0_C_5_io_in_lo = {IN_CHANX_N24232_70,IN_CHANX_N24222_30}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C37_N29303_O_0_C_5_io_in_hi = {IN_CHANY_N29399_37,IN_CHANX_N24270_50,IN_CHANX_N24260_10}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C45_N29311_O_0_C_5_io_in_lo = {IN_CHANX_N24208_52,IN_CHANX_N24198_12}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C45_N29311_O_0_C_5_io_in_hi = {IN_CHANY_N29401_45,IN_CHANX_N24254_72,IN_CHANX_N24244_32}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C53_N29319_O_0_C_5_io_in_lo = {IN_CHANX_N24228_54,IN_CHANX_N24218_14}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C53_N29319_O_0_C_5_io_in_hi = {IN_CHANY_N29403_53,IN_CHANX_N24276_74,IN_CHANX_N24266_34}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C61_N29327_O_0_C_5_io_in_lo = {IN_CHANX_N24240_16,IN_CHANX_N24204_36}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C61_N29327_O_0_C_5_io_in_hi = {IN_CHANY_N29405_61,IN_CHANX_N24256_76,IN_CHANX_N24250_56}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C69_N29335_O_0_C_5_io_in_lo = {IN_CHANX_N24262_18,IN_CHANX_N24224_38}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C69_N29335_O_0_C_5_io_in_hi = {IN_CHANY_N29407_69,IN_CHANX_N24278_78,IN_CHANX_N24272_58}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C77_N29367_O_0_C_5_io_in_lo = {IN_CHANX_N24210_60,IN_CHANX_N24200_20}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C77_N29367_O_0_C_5_io_in_hi = {IN_CHANY_N29409_77,IN_CHANX_N24246_40,IN_CHANX_N24236_0}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C4_N29390_O_0_C_5_io_in_hi = {IN_CHANY_N29270_4,IN_CHANX_N24246_40,IN_CHANX_N24236_0}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C12_N29392_O_0_C_5_io_in_hi = {IN_CHANY_N29278_12,IN_CHANX_N24278_78,IN_CHANX_N24272_58}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C20_N29394_O_0_C_5_io_in_hi = {IN_CHANY_N29286_20,IN_CHANX_N24256_76,IN_CHANX_N24250_56}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C28_N29396_O_0_C_5_io_in_hi = {IN_CHANY_N29294_28,IN_CHANX_N24276_74,IN_CHANX_N24266_34}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C36_N29398_O_0_C_5_io_in_hi = {IN_CHANY_N29302_36,IN_CHANX_N24254_72,IN_CHANX_N24244_32}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C44_N29400_O_0_C_5_io_in_hi = {IN_CHANY_N29310_44,IN_CHANX_N24270_50,IN_CHANX_N24260_10}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C52_N29402_O_0_C_5_io_in_hi = {IN_CHANY_N29318_52,IN_CHANX_N24248_48,IN_CHANX_N24238_8}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C60_N29404_O_0_C_5_io_in_hi = {IN_CHANY_N29326_60,IN_CHANX_N24274_66,IN_CHANX_N24264_26}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C68_N29406_O_0_C_5_io_in_hi = {IN_CHANY_N29334_68,IN_CHANX_N24252_64,IN_CHANX_N24242_24}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C76_N29408_O_0_C_5_io_in_hi = {IN_CHANY_N29366_76,IN_CHANX_N24268_42,IN_CHANX_N24258_2}; // @[TileFull.scala 183:11]
  IOBlock logicBlock ( // @[TileFull.scala 44:33]
    .IPIN_0(logicBlock_IPIN_0),
    .IPIN_2(logicBlock_IPIN_2),
    .IPIN_4(logicBlock_IPIN_4),
    .IPIN_6(logicBlock_IPIN_6),
    .IPIN_8(logicBlock_IPIN_8),
    .IPIN_10(logicBlock_IPIN_10),
    .IPIN_12(logicBlock_IPIN_12),
    .IPIN_14(logicBlock_IPIN_14),
    .IPIN_16(logicBlock_IPIN_16),
    .IPIN_18(logicBlock_IPIN_18),
    .IPIN_20(logicBlock_IPIN_20),
    .IPIN_22(logicBlock_IPIN_22),
    .IPIN_24(logicBlock_IPIN_24),
    .IPIN_26(logicBlock_IPIN_26),
    .IPIN_28(logicBlock_IPIN_28),
    .IPIN_30(logicBlock_IPIN_30),
    .IPIN_32(logicBlock_IPIN_32),
    .IPIN_34(logicBlock_IPIN_34),
    .IPIN_36(logicBlock_IPIN_36),
    .IPIN_38(logicBlock_IPIN_38),
    .IPIN_40(logicBlock_IPIN_40),
    .IPIN_42(logicBlock_IPIN_42),
    .IPIN_44(logicBlock_IPIN_44),
    .IPIN_46(logicBlock_IPIN_46),
    .IPIN_48(logicBlock_IPIN_48),
    .IPIN_50(logicBlock_IPIN_50),
    .IPIN_52(logicBlock_IPIN_52),
    .IPIN_54(logicBlock_IPIN_54),
    .IPIN_56(logicBlock_IPIN_56),
    .IPIN_58(logicBlock_IPIN_58),
    .IPIN_60(logicBlock_IPIN_60),
    .IPIN_62(logicBlock_IPIN_62),
    .OPIN_1(logicBlock_OPIN_1),
    .OPIN_3(logicBlock_OPIN_3),
    .OPIN_5(logicBlock_OPIN_5),
    .OPIN_7(logicBlock_OPIN_7),
    .OPIN_9(logicBlock_OPIN_9),
    .OPIN_11(logicBlock_OPIN_11),
    .OPIN_13(logicBlock_OPIN_13),
    .OPIN_15(logicBlock_OPIN_15),
    .OPIN_17(logicBlock_OPIN_17),
    .OPIN_19(logicBlock_OPIN_19),
    .OPIN_21(logicBlock_OPIN_21),
    .OPIN_23(logicBlock_OPIN_23),
    .OPIN_25(logicBlock_OPIN_25),
    .OPIN_27(logicBlock_OPIN_27),
    .OPIN_29(logicBlock_OPIN_29),
    .OPIN_31(logicBlock_OPIN_31),
    .OPIN_33(logicBlock_OPIN_33),
    .OPIN_35(logicBlock_OPIN_35),
    .OPIN_37(logicBlock_OPIN_37),
    .OPIN_39(logicBlock_OPIN_39),
    .OPIN_41(logicBlock_OPIN_41),
    .OPIN_43(logicBlock_OPIN_43),
    .OPIN_45(logicBlock_OPIN_45),
    .OPIN_47(logicBlock_OPIN_47),
    .OPIN_49(logicBlock_OPIN_49),
    .OPIN_51(logicBlock_OPIN_51),
    .OPIN_53(logicBlock_OPIN_53),
    .OPIN_55(logicBlock_OPIN_55),
    .OPIN_57(logicBlock_OPIN_57),
    .OPIN_59(logicBlock_OPIN_59),
    .OPIN_61(logicBlock_OPIN_61),
    .OPIN_63(logicBlock_OPIN_63),
    .clock(logicBlock_clock),
    .reset(logicBlock_reset),
    .ioPad_i(logicBlock_ioPad_i),
    .ioPad_o(logicBlock_ioPad_o),
    .configBits(logicBlock_configBits),
    .loopBreak(logicBlock_loopBreak),
    .gndLBouts(logicBlock_gndLBouts)
  );
  ScanConf_Tile_11_3_iotile configBlock ( // @[TileFull.scala 61:31]
    .clock(configBlock_clock),
    .ioBundle_confOut(configBlock_ioBundle_confOut),
    .ioBundle_scan_in(configBlock_ioBundle_scan_in),
    .ioBundle_scan_en(configBlock_ioBundle_scan_en),
    .ioBundle_scan_out(configBlock_ioBundle_scan_out)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN0_N22160 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN0_N22160_io_in),
    .io_config(CBMux_IPIN0_N22160_io_config),
    .io_out(CBMux_IPIN0_N22160_io_out),
    .io_loopBreak(CBMux_IPIN0_N22160_io_loopBreak),
    .io_cnstClk(CBMux_IPIN0_N22160_io_cnstClk),
    .io_arst(CBMux_IPIN0_N22160_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN2_N22162 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN2_N22162_io_in),
    .io_config(CBMux_IPIN2_N22162_io_config),
    .io_out(CBMux_IPIN2_N22162_io_out),
    .io_loopBreak(CBMux_IPIN2_N22162_io_loopBreak),
    .io_cnstClk(CBMux_IPIN2_N22162_io_cnstClk),
    .io_arst(CBMux_IPIN2_N22162_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN4_N22164 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN4_N22164_io_in),
    .io_config(CBMux_IPIN4_N22164_io_config),
    .io_out(CBMux_IPIN4_N22164_io_out),
    .io_loopBreak(CBMux_IPIN4_N22164_io_loopBreak),
    .io_cnstClk(CBMux_IPIN4_N22164_io_cnstClk),
    .io_arst(CBMux_IPIN4_N22164_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN6_N22166 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN6_N22166_io_in),
    .io_config(CBMux_IPIN6_N22166_io_config),
    .io_out(CBMux_IPIN6_N22166_io_out),
    .io_loopBreak(CBMux_IPIN6_N22166_io_loopBreak),
    .io_cnstClk(CBMux_IPIN6_N22166_io_cnstClk),
    .io_arst(CBMux_IPIN6_N22166_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN8_N22168 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN8_N22168_io_in),
    .io_config(CBMux_IPIN8_N22168_io_config),
    .io_out(CBMux_IPIN8_N22168_io_out),
    .io_loopBreak(CBMux_IPIN8_N22168_io_loopBreak),
    .io_cnstClk(CBMux_IPIN8_N22168_io_cnstClk),
    .io_arst(CBMux_IPIN8_N22168_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN10_N22170 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN10_N22170_io_in),
    .io_config(CBMux_IPIN10_N22170_io_config),
    .io_out(CBMux_IPIN10_N22170_io_out),
    .io_loopBreak(CBMux_IPIN10_N22170_io_loopBreak),
    .io_cnstClk(CBMux_IPIN10_N22170_io_cnstClk),
    .io_arst(CBMux_IPIN10_N22170_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN12_N22172 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN12_N22172_io_in),
    .io_config(CBMux_IPIN12_N22172_io_config),
    .io_out(CBMux_IPIN12_N22172_io_out),
    .io_loopBreak(CBMux_IPIN12_N22172_io_loopBreak),
    .io_cnstClk(CBMux_IPIN12_N22172_io_cnstClk),
    .io_arst(CBMux_IPIN12_N22172_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN14_N22174 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN14_N22174_io_in),
    .io_config(CBMux_IPIN14_N22174_io_config),
    .io_out(CBMux_IPIN14_N22174_io_out),
    .io_loopBreak(CBMux_IPIN14_N22174_io_loopBreak),
    .io_cnstClk(CBMux_IPIN14_N22174_io_cnstClk),
    .io_arst(CBMux_IPIN14_N22174_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN16_N22176 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN16_N22176_io_in),
    .io_config(CBMux_IPIN16_N22176_io_config),
    .io_out(CBMux_IPIN16_N22176_io_out),
    .io_loopBreak(CBMux_IPIN16_N22176_io_loopBreak),
    .io_cnstClk(CBMux_IPIN16_N22176_io_cnstClk),
    .io_arst(CBMux_IPIN16_N22176_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN18_N22178 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN18_N22178_io_in),
    .io_config(CBMux_IPIN18_N22178_io_config),
    .io_out(CBMux_IPIN18_N22178_io_out),
    .io_loopBreak(CBMux_IPIN18_N22178_io_loopBreak),
    .io_cnstClk(CBMux_IPIN18_N22178_io_cnstClk),
    .io_arst(CBMux_IPIN18_N22178_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN20_N22180 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN20_N22180_io_in),
    .io_config(CBMux_IPIN20_N22180_io_config),
    .io_out(CBMux_IPIN20_N22180_io_out),
    .io_loopBreak(CBMux_IPIN20_N22180_io_loopBreak),
    .io_cnstClk(CBMux_IPIN20_N22180_io_cnstClk),
    .io_arst(CBMux_IPIN20_N22180_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN22_N22182 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN22_N22182_io_in),
    .io_config(CBMux_IPIN22_N22182_io_config),
    .io_out(CBMux_IPIN22_N22182_io_out),
    .io_loopBreak(CBMux_IPIN22_N22182_io_loopBreak),
    .io_cnstClk(CBMux_IPIN22_N22182_io_cnstClk),
    .io_arst(CBMux_IPIN22_N22182_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN24_N22184 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN24_N22184_io_in),
    .io_config(CBMux_IPIN24_N22184_io_config),
    .io_out(CBMux_IPIN24_N22184_io_out),
    .io_loopBreak(CBMux_IPIN24_N22184_io_loopBreak),
    .io_cnstClk(CBMux_IPIN24_N22184_io_cnstClk),
    .io_arst(CBMux_IPIN24_N22184_io_arst)
  );
  MuxNInput_20_SCAOptCB CBMux_IPIN26_N22186 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN26_N22186_io_in),
    .io_config(CBMux_IPIN26_N22186_io_config),
    .io_out(CBMux_IPIN26_N22186_io_out),
    .io_loopBreak(CBMux_IPIN26_N22186_io_loopBreak),
    .io_cnstClk(CBMux_IPIN26_N22186_io_cnstClk),
    .io_arst(CBMux_IPIN26_N22186_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN28_N22188 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN28_N22188_io_in),
    .io_config(CBMux_IPIN28_N22188_io_config),
    .io_out(CBMux_IPIN28_N22188_io_out),
    .io_loopBreak(CBMux_IPIN28_N22188_io_loopBreak),
    .io_cnstClk(CBMux_IPIN28_N22188_io_cnstClk),
    .io_arst(CBMux_IPIN28_N22188_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN30_N22190 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN30_N22190_io_in),
    .io_config(CBMux_IPIN30_N22190_io_config),
    .io_out(CBMux_IPIN30_N22190_io_out),
    .io_loopBreak(CBMux_IPIN30_N22190_io_loopBreak),
    .io_cnstClk(CBMux_IPIN30_N22190_io_cnstClk),
    .io_arst(CBMux_IPIN30_N22190_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN32_N22192 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN32_N22192_io_in),
    .io_config(CBMux_IPIN32_N22192_io_config),
    .io_out(CBMux_IPIN32_N22192_io_out),
    .io_loopBreak(CBMux_IPIN32_N22192_io_loopBreak),
    .io_cnstClk(CBMux_IPIN32_N22192_io_cnstClk),
    .io_arst(CBMux_IPIN32_N22192_io_arst)
  );
  MuxNInput_20_SCAOptCB CBMux_IPIN34_N22194 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN34_N22194_io_in),
    .io_config(CBMux_IPIN34_N22194_io_config),
    .io_out(CBMux_IPIN34_N22194_io_out),
    .io_loopBreak(CBMux_IPIN34_N22194_io_loopBreak),
    .io_cnstClk(CBMux_IPIN34_N22194_io_cnstClk),
    .io_arst(CBMux_IPIN34_N22194_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN36_N22196 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN36_N22196_io_in),
    .io_config(CBMux_IPIN36_N22196_io_config),
    .io_out(CBMux_IPIN36_N22196_io_out),
    .io_loopBreak(CBMux_IPIN36_N22196_io_loopBreak),
    .io_cnstClk(CBMux_IPIN36_N22196_io_cnstClk),
    .io_arst(CBMux_IPIN36_N22196_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN38_N22198 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN38_N22198_io_in),
    .io_config(CBMux_IPIN38_N22198_io_config),
    .io_out(CBMux_IPIN38_N22198_io_out),
    .io_loopBreak(CBMux_IPIN38_N22198_io_loopBreak),
    .io_cnstClk(CBMux_IPIN38_N22198_io_cnstClk),
    .io_arst(CBMux_IPIN38_N22198_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN40_N22200 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN40_N22200_io_in),
    .io_config(CBMux_IPIN40_N22200_io_config),
    .io_out(CBMux_IPIN40_N22200_io_out),
    .io_loopBreak(CBMux_IPIN40_N22200_io_loopBreak),
    .io_cnstClk(CBMux_IPIN40_N22200_io_cnstClk),
    .io_arst(CBMux_IPIN40_N22200_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN42_N22202 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN42_N22202_io_in),
    .io_config(CBMux_IPIN42_N22202_io_config),
    .io_out(CBMux_IPIN42_N22202_io_out),
    .io_loopBreak(CBMux_IPIN42_N22202_io_loopBreak),
    .io_cnstClk(CBMux_IPIN42_N22202_io_cnstClk),
    .io_arst(CBMux_IPIN42_N22202_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN44_N22204 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN44_N22204_io_in),
    .io_config(CBMux_IPIN44_N22204_io_config),
    .io_out(CBMux_IPIN44_N22204_io_out),
    .io_loopBreak(CBMux_IPIN44_N22204_io_loopBreak),
    .io_cnstClk(CBMux_IPIN44_N22204_io_cnstClk),
    .io_arst(CBMux_IPIN44_N22204_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN46_N22206 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN46_N22206_io_in),
    .io_config(CBMux_IPIN46_N22206_io_config),
    .io_out(CBMux_IPIN46_N22206_io_out),
    .io_loopBreak(CBMux_IPIN46_N22206_io_loopBreak),
    .io_cnstClk(CBMux_IPIN46_N22206_io_cnstClk),
    .io_arst(CBMux_IPIN46_N22206_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN48_N22208 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN48_N22208_io_in),
    .io_config(CBMux_IPIN48_N22208_io_config),
    .io_out(CBMux_IPIN48_N22208_io_out),
    .io_loopBreak(CBMux_IPIN48_N22208_io_loopBreak),
    .io_cnstClk(CBMux_IPIN48_N22208_io_cnstClk),
    .io_arst(CBMux_IPIN48_N22208_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN50_N22210 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN50_N22210_io_in),
    .io_config(CBMux_IPIN50_N22210_io_config),
    .io_out(CBMux_IPIN50_N22210_io_out),
    .io_loopBreak(CBMux_IPIN50_N22210_io_loopBreak),
    .io_cnstClk(CBMux_IPIN50_N22210_io_cnstClk),
    .io_arst(CBMux_IPIN50_N22210_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN52_N22212 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN52_N22212_io_in),
    .io_config(CBMux_IPIN52_N22212_io_config),
    .io_out(CBMux_IPIN52_N22212_io_out),
    .io_loopBreak(CBMux_IPIN52_N22212_io_loopBreak),
    .io_cnstClk(CBMux_IPIN52_N22212_io_cnstClk),
    .io_arst(CBMux_IPIN52_N22212_io_arst)
  );
  MuxNInput_16_SCAOptCB CBMux_IPIN54_N22214 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN54_N22214_io_in),
    .io_config(CBMux_IPIN54_N22214_io_config),
    .io_out(CBMux_IPIN54_N22214_io_out),
    .io_loopBreak(CBMux_IPIN54_N22214_io_loopBreak),
    .io_cnstClk(CBMux_IPIN54_N22214_io_cnstClk),
    .io_arst(CBMux_IPIN54_N22214_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN56_N22216 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN56_N22216_io_in),
    .io_config(CBMux_IPIN56_N22216_io_config),
    .io_out(CBMux_IPIN56_N22216_io_out),
    .io_loopBreak(CBMux_IPIN56_N22216_io_loopBreak),
    .io_cnstClk(CBMux_IPIN56_N22216_io_cnstClk),
    .io_arst(CBMux_IPIN56_N22216_io_arst)
  );
  MuxNInput_20_SCAOptCB CBMux_IPIN58_N22218 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN58_N22218_io_in),
    .io_config(CBMux_IPIN58_N22218_io_config),
    .io_out(CBMux_IPIN58_N22218_io_out),
    .io_loopBreak(CBMux_IPIN58_N22218_io_loopBreak),
    .io_cnstClk(CBMux_IPIN58_N22218_io_cnstClk),
    .io_arst(CBMux_IPIN58_N22218_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN60_N22220 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN60_N22220_io_in),
    .io_config(CBMux_IPIN60_N22220_io_config),
    .io_out(CBMux_IPIN60_N22220_io_out),
    .io_loopBreak(CBMux_IPIN60_N22220_io_loopBreak),
    .io_cnstClk(CBMux_IPIN60_N22220_io_cnstClk),
    .io_arst(CBMux_IPIN60_N22220_io_arst)
  );
  MuxNInput_18_SCAOptCB CBMux_IPIN62_N22222 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN62_N22222_io_in),
    .io_config(CBMux_IPIN62_N22222_io_config),
    .io_out(CBMux_IPIN62_N22222_io_out),
    .io_loopBreak(CBMux_IPIN62_N22222_io_loopBreak),
    .io_cnstClk(CBMux_IPIN62_N22222_io_cnstClk),
    .io_arst(CBMux_IPIN62_N22222_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C5_N24197_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C5_N24197_O_7_C_1_io_in),
    .io_config(SBMux_C5_N24197_O_7_C_1_io_config),
    .io_out(SBMux_C5_N24197_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C5_N24197_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C5_N24197_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C5_N24197_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C5_N24197_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C13_N24199_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C13_N24199_O_7_C_1_io_in),
    .io_config(SBMux_C13_N24199_O_7_C_1_io_config),
    .io_out(SBMux_C13_N24199_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C13_N24199_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C13_N24199_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C13_N24199_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C13_N24199_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C21_N24201_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C21_N24201_O_7_C_1_io_in),
    .io_config(SBMux_C21_N24201_O_7_C_1_io_config),
    .io_out(SBMux_C21_N24201_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C21_N24201_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C21_N24201_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C21_N24201_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C21_N24201_O_7_C_1_io_arst)
  );
  MuxNInput_O6_C1_SCAOptSB SBMux_C29_N24203_O_6_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C29_N24203_O_6_C_1_io_in),
    .io_config(SBMux_C29_N24203_O_6_C_1_io_config),
    .io_out(SBMux_C29_N24203_O_6_C_1_io_out),
    .io_loopBreak(SBMux_C29_N24203_O_6_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C29_N24203_O_6_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C29_N24203_O_6_C_1_io_cnstClk),
    .io_arst(SBMux_C29_N24203_O_6_C_1_io_arst)
  );
  MuxNInput_O6_C2_SCAOptSB SBMux_C37_N24205_O_6_C_2 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C37_N24205_O_6_C_2_io_in),
    .io_config(SBMux_C37_N24205_O_6_C_2_io_config),
    .io_out(SBMux_C37_N24205_O_6_C_2_io_out),
    .io_loopBreak(SBMux_C37_N24205_O_6_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C37_N24205_O_6_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C37_N24205_O_6_C_2_io_cnstClk),
    .io_arst(SBMux_C37_N24205_O_6_C_2_io_arst)
  );
  MuxNInput_O7_C2_SCAOptSB SBMux_C45_N24207_O_7_C_2 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C45_N24207_O_7_C_2_io_in),
    .io_config(SBMux_C45_N24207_O_7_C_2_io_config),
    .io_out(SBMux_C45_N24207_O_7_C_2_io_out),
    .io_loopBreak(SBMux_C45_N24207_O_7_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C45_N24207_O_7_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C45_N24207_O_7_C_2_io_cnstClk),
    .io_arst(SBMux_C45_N24207_O_7_C_2_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C53_N24209_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C53_N24209_O_7_C_1_io_in),
    .io_config(SBMux_C53_N24209_O_7_C_1_io_config),
    .io_out(SBMux_C53_N24209_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C53_N24209_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C53_N24209_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C53_N24209_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C53_N24209_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C61_N24211_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C61_N24211_O_7_C_1_io_in),
    .io_config(SBMux_C61_N24211_O_7_C_1_io_config),
    .io_out(SBMux_C61_N24211_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C61_N24211_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C61_N24211_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C61_N24211_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C61_N24211_O_7_C_1_io_arst)
  );
  MuxNInput_O6_C1_SCAOptSB SBMux_C69_N24213_O_6_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C69_N24213_O_6_C_1_io_in),
    .io_config(SBMux_C69_N24213_O_6_C_1_io_config),
    .io_out(SBMux_C69_N24213_O_6_C_1_io_out),
    .io_loopBreak(SBMux_C69_N24213_O_6_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C69_N24213_O_6_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C69_N24213_O_6_C_1_io_cnstClk),
    .io_arst(SBMux_C69_N24213_O_6_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C7_N24217_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C7_N24217_O_7_C_1_io_in),
    .io_config(SBMux_C7_N24217_O_7_C_1_io_config),
    .io_out(SBMux_C7_N24217_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C7_N24217_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C7_N24217_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C7_N24217_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C7_N24217_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C15_N24219_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C15_N24219_O_7_C_1_io_in),
    .io_config(SBMux_C15_N24219_O_7_C_1_io_config),
    .io_out(SBMux_C15_N24219_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C15_N24219_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C15_N24219_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C15_N24219_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C15_N24219_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C23_N24221_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C23_N24221_O_7_C_1_io_in),
    .io_config(SBMux_C23_N24221_O_7_C_1_io_config),
    .io_out(SBMux_C23_N24221_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C23_N24221_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C23_N24221_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C23_N24221_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C23_N24221_O_7_C_1_io_arst)
  );
  MuxNInput_O6_C1_SCAOptSB SBMux_C31_N24223_O_6_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C31_N24223_O_6_C_1_io_in),
    .io_config(SBMux_C31_N24223_O_6_C_1_io_config),
    .io_out(SBMux_C31_N24223_O_6_C_1_io_out),
    .io_loopBreak(SBMux_C31_N24223_O_6_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C31_N24223_O_6_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C31_N24223_O_6_C_1_io_cnstClk),
    .io_arst(SBMux_C31_N24223_O_6_C_1_io_arst)
  );
  MuxNInput_O7_C2_SCAOptSB SBMux_C39_N24225_O_7_C_2 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C39_N24225_O_7_C_2_io_in),
    .io_config(SBMux_C39_N24225_O_7_C_2_io_config),
    .io_out(SBMux_C39_N24225_O_7_C_2_io_out),
    .io_loopBreak(SBMux_C39_N24225_O_7_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C39_N24225_O_7_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C39_N24225_O_7_C_2_io_cnstClk),
    .io_arst(SBMux_C39_N24225_O_7_C_2_io_arst)
  );
  MuxNInput_O7_C2_SCAOptSB SBMux_C47_N24227_O_7_C_2 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C47_N24227_O_7_C_2_io_in),
    .io_config(SBMux_C47_N24227_O_7_C_2_io_config),
    .io_out(SBMux_C47_N24227_O_7_C_2_io_out),
    .io_loopBreak(SBMux_C47_N24227_O_7_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C47_N24227_O_7_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C47_N24227_O_7_C_2_io_cnstClk),
    .io_arst(SBMux_C47_N24227_O_7_C_2_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C55_N24229_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C55_N24229_O_7_C_1_io_in),
    .io_config(SBMux_C55_N24229_O_7_C_1_io_config),
    .io_out(SBMux_C55_N24229_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C55_N24229_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C55_N24229_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C55_N24229_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C55_N24229_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C63_N24231_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C63_N24231_O_7_C_1_io_in),
    .io_config(SBMux_C63_N24231_O_7_C_1_io_config),
    .io_out(SBMux_C63_N24231_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C63_N24231_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C63_N24231_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C63_N24231_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C63_N24231_O_7_C_1_io_arst)
  );
  MuxNInput_O6_C1_SCAOptSB SBMux_C71_N24233_O_6_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C71_N24233_O_6_C_1_io_in),
    .io_config(SBMux_C71_N24233_O_6_C_1_io_config),
    .io_out(SBMux_C71_N24233_O_6_C_1_io_out),
    .io_loopBreak(SBMux_C71_N24233_O_6_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C71_N24233_O_6_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C71_N24233_O_6_C_1_io_cnstClk),
    .io_arst(SBMux_C71_N24233_O_6_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C1_N24237_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C1_N24237_O_7_C_1_io_in),
    .io_config(SBMux_C1_N24237_O_7_C_1_io_config),
    .io_out(SBMux_C1_N24237_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C1_N24237_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C1_N24237_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C1_N24237_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C1_N24237_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C9_N24239_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C9_N24239_O_7_C_1_io_in),
    .io_config(SBMux_C9_N24239_O_7_C_1_io_config),
    .io_out(SBMux_C9_N24239_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C9_N24239_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C9_N24239_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C9_N24239_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C9_N24239_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C17_N24241_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C17_N24241_O_7_C_1_io_in),
    .io_config(SBMux_C17_N24241_O_7_C_1_io_config),
    .io_out(SBMux_C17_N24241_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C17_N24241_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C17_N24241_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C17_N24241_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C17_N24241_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C25_N24243_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C25_N24243_O_7_C_1_io_in),
    .io_config(SBMux_C25_N24243_O_7_C_1_io_config),
    .io_out(SBMux_C25_N24243_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C25_N24243_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C25_N24243_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C25_N24243_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C25_N24243_O_7_C_1_io_arst)
  );
  MuxNInput_O6_C1_SCAOptSB SBMux_C33_N24245_O_6_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C33_N24245_O_6_C_1_io_in),
    .io_config(SBMux_C33_N24245_O_6_C_1_io_config),
    .io_out(SBMux_C33_N24245_O_6_C_1_io_out),
    .io_loopBreak(SBMux_C33_N24245_O_6_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C33_N24245_O_6_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C33_N24245_O_6_C_1_io_cnstClk),
    .io_arst(SBMux_C33_N24245_O_6_C_1_io_arst)
  );
  MuxNInput_O7_C2_SCAOptSB SBMux_C41_N24247_O_7_C_2 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C41_N24247_O_7_C_2_io_in),
    .io_config(SBMux_C41_N24247_O_7_C_2_io_config),
    .io_out(SBMux_C41_N24247_O_7_C_2_io_out),
    .io_loopBreak(SBMux_C41_N24247_O_7_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C41_N24247_O_7_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C41_N24247_O_7_C_2_io_cnstClk),
    .io_arst(SBMux_C41_N24247_O_7_C_2_io_arst)
  );
  MuxNInput_O7_C2_SCAOptSB SBMux_C49_N24249_O_7_C_2 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C49_N24249_O_7_C_2_io_in),
    .io_config(SBMux_C49_N24249_O_7_C_2_io_config),
    .io_out(SBMux_C49_N24249_O_7_C_2_io_out),
    .io_loopBreak(SBMux_C49_N24249_O_7_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C49_N24249_O_7_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C49_N24249_O_7_C_2_io_cnstClk),
    .io_arst(SBMux_C49_N24249_O_7_C_2_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C57_N24251_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C57_N24251_O_7_C_1_io_in),
    .io_config(SBMux_C57_N24251_O_7_C_1_io_config),
    .io_out(SBMux_C57_N24251_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C57_N24251_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C57_N24251_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C57_N24251_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C57_N24251_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C65_N24253_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C65_N24253_O_7_C_1_io_in),
    .io_config(SBMux_C65_N24253_O_7_C_1_io_config),
    .io_out(SBMux_C65_N24253_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C65_N24253_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C65_N24253_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C65_N24253_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C65_N24253_O_7_C_1_io_arst)
  );
  MuxNInput_O6_C1_SCAOptSB SBMux_C73_N24255_O_6_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C73_N24255_O_6_C_1_io_in),
    .io_config(SBMux_C73_N24255_O_6_C_1_io_config),
    .io_out(SBMux_C73_N24255_O_6_C_1_io_out),
    .io_loopBreak(SBMux_C73_N24255_O_6_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C73_N24255_O_6_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C73_N24255_O_6_C_1_io_cnstClk),
    .io_arst(SBMux_C73_N24255_O_6_C_1_io_arst)
  );
  MuxNInput_O16_C1_SCAOptSB SBMux_C77_N24257_O_16_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C77_N24257_O_16_C_1_io_in),
    .io_config(SBMux_C77_N24257_O_16_C_1_io_config),
    .io_out(SBMux_C77_N24257_O_16_C_1_io_out),
    .io_loopBreak(SBMux_C77_N24257_O_16_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C77_N24257_O_16_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C77_N24257_O_16_C_1_io_cnstClk),
    .io_arst(SBMux_C77_N24257_O_16_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C3_N24259_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C3_N24259_O_7_C_1_io_in),
    .io_config(SBMux_C3_N24259_O_7_C_1_io_config),
    .io_out(SBMux_C3_N24259_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C3_N24259_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C3_N24259_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C3_N24259_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C3_N24259_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C11_N24261_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C11_N24261_O_7_C_1_io_in),
    .io_config(SBMux_C11_N24261_O_7_C_1_io_config),
    .io_out(SBMux_C11_N24261_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C11_N24261_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C11_N24261_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C11_N24261_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C11_N24261_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C19_N24263_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C19_N24263_O_7_C_1_io_in),
    .io_config(SBMux_C19_N24263_O_7_C_1_io_config),
    .io_out(SBMux_C19_N24263_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C19_N24263_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C19_N24263_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C19_N24263_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C19_N24263_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C27_N24265_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C27_N24265_O_7_C_1_io_in),
    .io_config(SBMux_C27_N24265_O_7_C_1_io_config),
    .io_out(SBMux_C27_N24265_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C27_N24265_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C27_N24265_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C27_N24265_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C27_N24265_O_7_C_1_io_arst)
  );
  MuxNInput_O6_C2_SCAOptSB SBMux_C35_N24267_O_6_C_2 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C35_N24267_O_6_C_2_io_in),
    .io_config(SBMux_C35_N24267_O_6_C_2_io_config),
    .io_out(SBMux_C35_N24267_O_6_C_2_io_out),
    .io_loopBreak(SBMux_C35_N24267_O_6_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C35_N24267_O_6_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C35_N24267_O_6_C_2_io_cnstClk),
    .io_arst(SBMux_C35_N24267_O_6_C_2_io_arst)
  );
  MuxNInput_O7_C2_SCAOptSB SBMux_C43_N24269_O_7_C_2 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C43_N24269_O_7_C_2_io_in),
    .io_config(SBMux_C43_N24269_O_7_C_2_io_config),
    .io_out(SBMux_C43_N24269_O_7_C_2_io_out),
    .io_loopBreak(SBMux_C43_N24269_O_7_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C43_N24269_O_7_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C43_N24269_O_7_C_2_io_cnstClk),
    .io_arst(SBMux_C43_N24269_O_7_C_2_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C51_N24271_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C51_N24271_O_7_C_1_io_in),
    .io_config(SBMux_C51_N24271_O_7_C_1_io_config),
    .io_out(SBMux_C51_N24271_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C51_N24271_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C51_N24271_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C51_N24271_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C51_N24271_O_7_C_1_io_arst)
  );
  MuxNInput_O7_C1_SCAOptSB SBMux_C59_N24273_O_7_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C59_N24273_O_7_C_1_io_in),
    .io_config(SBMux_C59_N24273_O_7_C_1_io_config),
    .io_out(SBMux_C59_N24273_O_7_C_1_io_out),
    .io_loopBreak(SBMux_C59_N24273_O_7_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C59_N24273_O_7_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C59_N24273_O_7_C_1_io_cnstClk),
    .io_arst(SBMux_C59_N24273_O_7_C_1_io_arst)
  );
  MuxNInput_O6_C1_SCAOptSB SBMux_C67_N24275_O_6_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C67_N24275_O_6_C_1_io_in),
    .io_config(SBMux_C67_N24275_O_6_C_1_io_config),
    .io_out(SBMux_C67_N24275_O_6_C_1_io_out),
    .io_loopBreak(SBMux_C67_N24275_O_6_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C67_N24275_O_6_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C67_N24275_O_6_C_1_io_cnstClk),
    .io_arst(SBMux_C67_N24275_O_6_C_1_io_arst)
  );
  MuxNInput_O6_C1_SCAOptSB SBMux_C75_N24277_O_6_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C75_N24277_O_6_C_1_io_in),
    .io_config(SBMux_C75_N24277_O_6_C_1_io_config),
    .io_out(SBMux_C75_N24277_O_6_C_1_io_out),
    .io_loopBreak(SBMux_C75_N24277_O_6_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C75_N24277_O_6_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C75_N24277_O_6_C_1_io_cnstClk),
    .io_arst(SBMux_C75_N24277_O_6_C_1_io_arst)
  );
  MuxNInput_O16_C1_SCAOptSB SBMux_C79_N24279_O_16_C_1 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C79_N24279_O_16_C_1_io_in),
    .io_config(SBMux_C79_N24279_O_16_C_1_io_config),
    .io_out(SBMux_C79_N24279_O_16_C_1_io_out),
    .io_loopBreak(SBMux_C79_N24279_O_16_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C79_N24279_O_16_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C79_N24279_O_16_C_1_io_cnstClk),
    .io_arst(SBMux_C79_N24279_O_16_C_1_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C5_N29271_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C5_N29271_O_0_C_5_io_in),
    .io_config(SBMux_C5_N29271_O_0_C_5_io_config),
    .io_out(SBMux_C5_N29271_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C5_N29271_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C5_N29271_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C5_N29271_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C5_N29271_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C13_N29279_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C13_N29279_O_0_C_5_io_in),
    .io_config(SBMux_C13_N29279_O_0_C_5_io_config),
    .io_out(SBMux_C13_N29279_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C13_N29279_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C13_N29279_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C13_N29279_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C13_N29279_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C21_N29287_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C21_N29287_O_0_C_5_io_in),
    .io_config(SBMux_C21_N29287_O_0_C_5_io_config),
    .io_out(SBMux_C21_N29287_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C21_N29287_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C21_N29287_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C21_N29287_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C21_N29287_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C29_N29295_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C29_N29295_O_0_C_5_io_in),
    .io_config(SBMux_C29_N29295_O_0_C_5_io_config),
    .io_out(SBMux_C29_N29295_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C29_N29295_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C29_N29295_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C29_N29295_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C29_N29295_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C37_N29303_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C37_N29303_O_0_C_5_io_in),
    .io_config(SBMux_C37_N29303_O_0_C_5_io_config),
    .io_out(SBMux_C37_N29303_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C37_N29303_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C37_N29303_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C37_N29303_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C37_N29303_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C45_N29311_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C45_N29311_O_0_C_5_io_in),
    .io_config(SBMux_C45_N29311_O_0_C_5_io_config),
    .io_out(SBMux_C45_N29311_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C45_N29311_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C45_N29311_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C45_N29311_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C45_N29311_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C53_N29319_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C53_N29319_O_0_C_5_io_in),
    .io_config(SBMux_C53_N29319_O_0_C_5_io_config),
    .io_out(SBMux_C53_N29319_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C53_N29319_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C53_N29319_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C53_N29319_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C53_N29319_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C61_N29327_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C61_N29327_O_0_C_5_io_in),
    .io_config(SBMux_C61_N29327_O_0_C_5_io_config),
    .io_out(SBMux_C61_N29327_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C61_N29327_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C61_N29327_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C61_N29327_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C61_N29327_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C69_N29335_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C69_N29335_O_0_C_5_io_in),
    .io_config(SBMux_C69_N29335_O_0_C_5_io_config),
    .io_out(SBMux_C69_N29335_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C69_N29335_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C69_N29335_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C69_N29335_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C69_N29335_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C77_N29367_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C77_N29367_O_0_C_5_io_in),
    .io_config(SBMux_C77_N29367_O_0_C_5_io_config),
    .io_out(SBMux_C77_N29367_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C77_N29367_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C77_N29367_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C77_N29367_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C77_N29367_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C4_N29390_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C4_N29390_O_0_C_5_io_in),
    .io_config(SBMux_C4_N29390_O_0_C_5_io_config),
    .io_out(SBMux_C4_N29390_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C4_N29390_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C4_N29390_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C4_N29390_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C4_N29390_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C12_N29392_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C12_N29392_O_0_C_5_io_in),
    .io_config(SBMux_C12_N29392_O_0_C_5_io_config),
    .io_out(SBMux_C12_N29392_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C12_N29392_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C12_N29392_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C12_N29392_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C12_N29392_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C20_N29394_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C20_N29394_O_0_C_5_io_in),
    .io_config(SBMux_C20_N29394_O_0_C_5_io_config),
    .io_out(SBMux_C20_N29394_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C20_N29394_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C20_N29394_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C20_N29394_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C20_N29394_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C28_N29396_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C28_N29396_O_0_C_5_io_in),
    .io_config(SBMux_C28_N29396_O_0_C_5_io_config),
    .io_out(SBMux_C28_N29396_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C28_N29396_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C28_N29396_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C28_N29396_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C28_N29396_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C36_N29398_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C36_N29398_O_0_C_5_io_in),
    .io_config(SBMux_C36_N29398_O_0_C_5_io_config),
    .io_out(SBMux_C36_N29398_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C36_N29398_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C36_N29398_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C36_N29398_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C36_N29398_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C44_N29400_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C44_N29400_O_0_C_5_io_in),
    .io_config(SBMux_C44_N29400_O_0_C_5_io_config),
    .io_out(SBMux_C44_N29400_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C44_N29400_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C44_N29400_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C44_N29400_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C44_N29400_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C52_N29402_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C52_N29402_O_0_C_5_io_in),
    .io_config(SBMux_C52_N29402_O_0_C_5_io_config),
    .io_out(SBMux_C52_N29402_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C52_N29402_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C52_N29402_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C52_N29402_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C52_N29402_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C60_N29404_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C60_N29404_O_0_C_5_io_in),
    .io_config(SBMux_C60_N29404_O_0_C_5_io_config),
    .io_out(SBMux_C60_N29404_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C60_N29404_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C60_N29404_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C60_N29404_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C60_N29404_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C68_N29406_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C68_N29406_O_0_C_5_io_in),
    .io_config(SBMux_C68_N29406_O_0_C_5_io_config),
    .io_out(SBMux_C68_N29406_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C68_N29406_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C68_N29406_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C68_N29406_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C68_N29406_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C76_N29408_O_0_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C76_N29408_O_0_C_5_io_in),
    .io_config(SBMux_C76_N29408_O_0_C_5_io_config),
    .io_out(SBMux_C76_N29408_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C76_N29408_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C76_N29408_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C76_N29408_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C76_N29408_O_0_C_5_io_arst)
  );
  assign OUT_OPIN_N22211_51 = logicBlock_OPIN_51; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N29400_44 = SBMux_C44_N29400_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24229_55 = SBMux_C55_N24229_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24239_9 = SBMux_C9_N24239_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24269_43 = SBMux_C43_N24269_O_7_C_2_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29398_36 = SBMux_C36_N29398_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24237_1 = SBMux_C1_N24237_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24199_13 = SBMux_C13_N24199_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24211_61 = SBMux_C61_N24211_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22223_63 = logicBlock_OPIN_63; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24241_17 = SBMux_C17_N24241_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24213_69 = SBMux_C69_N24213_O_6_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24279_79 = SBMux_C79_N24279_O_16_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22193_33 = logicBlock_OPIN_33; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24207_45 = SBMux_C45_N24207_O_7_C_2_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22185_25 = logicBlock_OPIN_25; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24233_71 = SBMux_C71_N24233_O_6_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24221_23 = SBMux_C23_N24221_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24271_51 = SBMux_C51_N24271_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22187_27 = logicBlock_OPIN_27; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24245_33 = SBMux_C33_N24245_O_6_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24265_27 = SBMux_C27_N24265_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29390_4 = SBMux_C4_N29390_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29319_53 = SBMux_C53_N29319_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24209_53 = SBMux_C53_N24209_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24217_7 = SBMux_C7_N24217_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24273_59 = SBMux_C59_N24273_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29408_76 = SBMux_C76_N29408_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29287_21 = SBMux_C21_N29287_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24197_5 = SBMux_C5_N24197_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24267_35 = SBMux_C35_N24267_O_6_C_2_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24203_29 = SBMux_C29_N24203_O_6_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22183_23 = logicBlock_OPIN_23; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N29271_5 = SBMux_C5_N29271_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29406_68 = SBMux_C68_N29406_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24219_15 = SBMux_C15_N24219_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22161_1 = logicBlock_OPIN_1; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24201_21 = SBMux_C21_N24201_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22215_55 = logicBlock_OPIN_55; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24253_65 = SBMux_C65_N24253_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29295_29 = SBMux_C29_N29295_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22175_15 = logicBlock_OPIN_15; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22217_57 = logicBlock_OPIN_57; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22213_53 = logicBlock_OPIN_53; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N29303_37 = SBMux_C37_N29303_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29311_45 = SBMux_C45_N29311_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22177_17 = logicBlock_OPIN_17; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N29392_12 = SBMux_C12_N29392_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24205_37 = SBMux_C37_N24205_O_6_C_2_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24247_41 = SBMux_C41_N24247_O_7_C_2_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22163_3 = logicBlock_OPIN_3; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22165_5 = logicBlock_OPIN_5; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22189_29 = logicBlock_OPIN_29; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24255_73 = SBMux_C73_N24255_O_6_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24263_19 = SBMux_C19_N24263_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22169_9 = logicBlock_OPIN_9; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22207_47 = logicBlock_OPIN_47; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22201_41 = logicBlock_OPIN_41; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22205_45 = logicBlock_OPIN_45; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24251_57 = SBMux_C57_N24251_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22219_59 = logicBlock_OPIN_59; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N29402_52 = SBMux_C52_N29402_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29367_77 = SBMux_C77_N29367_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29394_20 = SBMux_C20_N29394_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24259_3 = SBMux_C3_N24259_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22221_61 = logicBlock_OPIN_61; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24223_31 = SBMux_C31_N24223_O_6_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24231_63 = SBMux_C63_N24231_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22181_21 = logicBlock_OPIN_21; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N29404_60 = SBMux_C60_N29404_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29327_61 = SBMux_C61_N29327_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22171_11 = logicBlock_OPIN_11; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24261_11 = SBMux_C11_N24261_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22195_35 = logicBlock_OPIN_35; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22179_19 = logicBlock_OPIN_19; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24275_67 = SBMux_C67_N24275_O_6_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N29396_28 = SBMux_C28_N29396_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24243_25 = SBMux_C25_N24243_O_7_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22167_7 = logicBlock_OPIN_7; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22197_37 = logicBlock_OPIN_37; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22209_49 = logicBlock_OPIN_49; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N29279_13 = SBMux_C13_N29279_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24277_75 = SBMux_C75_N24277_O_6_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22199_39 = logicBlock_OPIN_39; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24249_49 = SBMux_C49_N24249_O_7_C_2_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22203_43 = logicBlock_OPIN_43; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N22173_13 = logicBlock_OPIN_13; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N29335_69 = SBMux_C69_N29335_O_0_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24227_47 = SBMux_C47_N24227_O_7_C_2_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24257_77 = SBMux_C77_N24257_O_16_C_1_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24225_39 = SBMux_C39_N24225_O_7_C_2_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N22191_31 = logicBlock_OPIN_31; // @[TileFull.scala 196:12]
  assign ioConf_confOut = configBlock_ioBundle_confOut[417:0]; // @[TileFull.scala 73:12]
  assign ioConf_scan_out = configBlock_ioBundle_scan_out; // @[TileFull.scala 73:12]
  assign ioPad_o = logicBlock_ioPad_o; // @[TileFull.scala 202:15]
  assign logicBlock_IPIN_0 = CBMux_IPIN0_N22160_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_2 = CBMux_IPIN2_N22162_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_4 = CBMux_IPIN4_N22164_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_6 = CBMux_IPIN6_N22166_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_8 = CBMux_IPIN8_N22168_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_10 = CBMux_IPIN10_N22170_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_12 = CBMux_IPIN12_N22172_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_14 = CBMux_IPIN14_N22174_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_16 = CBMux_IPIN16_N22176_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_18 = CBMux_IPIN18_N22178_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_20 = CBMux_IPIN20_N22180_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_22 = CBMux_IPIN22_N22182_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_24 = CBMux_IPIN24_N22184_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_26 = CBMux_IPIN26_N22186_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_28 = CBMux_IPIN28_N22188_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_30 = CBMux_IPIN30_N22190_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_32 = CBMux_IPIN32_N22192_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_34 = CBMux_IPIN34_N22194_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_36 = CBMux_IPIN36_N22196_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_38 = CBMux_IPIN38_N22198_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_40 = CBMux_IPIN40_N22200_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_42 = CBMux_IPIN42_N22202_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_44 = CBMux_IPIN44_N22204_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_46 = CBMux_IPIN46_N22206_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_48 = CBMux_IPIN48_N22208_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_50 = CBMux_IPIN50_N22210_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_52 = CBMux_IPIN52_N22212_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_54 = CBMux_IPIN54_N22214_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_56 = CBMux_IPIN56_N22216_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_58 = CBMux_IPIN58_N22218_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_60 = CBMux_IPIN60_N22220_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_62 = CBMux_IPIN62_N22222_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_clock = clock; // @[TileFull.scala 192:26]
  assign logicBlock_reset = reset; // @[TileFull.scala 193:26]
  assign logicBlock_ioPad_i = ioPad_i; // @[TileFull.scala 202:15]
  assign logicBlock_configBits = configBlock_ioBundle_confOut[15:0]; // @[TileFull.scala 191:31]
  assign logicBlock_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 190:30]
  assign logicBlock_gndLBouts = ctrlSignals_gndBlkOuts; // @[TileFull.scala 189:30]
  assign configBlock_clock = ctrlSignals_confClock; // @[TileFull.scala 74:27]
  assign configBlock_ioBundle_scan_in = ioConf_scan_in; // @[TileFull.scala 73:12]
  assign configBlock_ioBundle_scan_en = ioConf_scan_en; // @[TileFull.scala 73:12]
  assign CBMux_IPIN0_N22160_io_in = {CBMux_IPIN0_N22160_io_in_hi,CBMux_IPIN0_N22160_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN0_N22160_io_config = configBlock_ioBundle_confOut[20:16]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN0_N22160_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN0_N22160_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN0_N22160_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN2_N22162_io_in = {CBMux_IPIN2_N22162_io_in_hi,CBMux_IPIN2_N22162_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN2_N22162_io_config = configBlock_ioBundle_confOut[25:21]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN2_N22162_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN2_N22162_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN2_N22162_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN4_N22164_io_in = {CBMux_IPIN4_N22164_io_in_hi,CBMux_IPIN4_N22164_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN4_N22164_io_config = configBlock_ioBundle_confOut[30:26]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN4_N22164_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN4_N22164_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN4_N22164_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN6_N22166_io_in = {CBMux_IPIN6_N22166_io_in_hi,CBMux_IPIN6_N22166_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN6_N22166_io_config = configBlock_ioBundle_confOut[35:31]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN6_N22166_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN6_N22166_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN6_N22166_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN8_N22168_io_in = {CBMux_IPIN8_N22168_io_in_hi,CBMux_IPIN8_N22168_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN8_N22168_io_config = configBlock_ioBundle_confOut[40:36]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN8_N22168_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN8_N22168_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN8_N22168_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN10_N22170_io_in = {CBMux_IPIN10_N22170_io_in_hi,CBMux_IPIN10_N22170_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN10_N22170_io_config = configBlock_ioBundle_confOut[45:41]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN10_N22170_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN10_N22170_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN10_N22170_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN12_N22172_io_in = {CBMux_IPIN12_N22172_io_in_hi,CBMux_IPIN12_N22172_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN12_N22172_io_config = configBlock_ioBundle_confOut[50:46]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN12_N22172_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN12_N22172_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN12_N22172_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN14_N22174_io_in = {CBMux_IPIN14_N22174_io_in_hi,CBMux_IPIN14_N22174_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN14_N22174_io_config = configBlock_ioBundle_confOut[55:51]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN14_N22174_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN14_N22174_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN14_N22174_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN16_N22176_io_in = {CBMux_IPIN16_N22176_io_in_hi,CBMux_IPIN16_N22176_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN16_N22176_io_config = configBlock_ioBundle_confOut[60:56]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN16_N22176_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN16_N22176_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN16_N22176_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN18_N22178_io_in = {CBMux_IPIN18_N22178_io_in_hi,CBMux_IPIN18_N22178_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN18_N22178_io_config = configBlock_ioBundle_confOut[65:61]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN18_N22178_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN18_N22178_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN18_N22178_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN20_N22180_io_in = {CBMux_IPIN20_N22180_io_in_hi,CBMux_IPIN20_N22180_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN20_N22180_io_config = configBlock_ioBundle_confOut[70:66]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN20_N22180_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN20_N22180_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN20_N22180_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN22_N22182_io_in = {CBMux_IPIN22_N22182_io_in_hi,CBMux_IPIN22_N22182_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN22_N22182_io_config = configBlock_ioBundle_confOut[75:71]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN22_N22182_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN22_N22182_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN22_N22182_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN24_N22184_io_in = {CBMux_IPIN24_N22184_io_in_hi,CBMux_IPIN24_N22184_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN24_N22184_io_config = configBlock_ioBundle_confOut[80:76]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN24_N22184_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN24_N22184_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN24_N22184_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN26_N22186_io_in = {CBMux_IPIN26_N22186_io_in_hi,CBMux_IPIN26_N22186_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN26_N22186_io_config = configBlock_ioBundle_confOut[85:81]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN26_N22186_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN26_N22186_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN26_N22186_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN28_N22188_io_in = {CBMux_IPIN20_N22180_io_in_hi,CBMux_IPIN28_N22188_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN28_N22188_io_config = configBlock_ioBundle_confOut[90:86]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN28_N22188_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN28_N22188_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN28_N22188_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN30_N22190_io_in = {CBMux_IPIN30_N22190_io_in_hi,CBMux_IPIN30_N22190_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN30_N22190_io_config = configBlock_ioBundle_confOut[95:91]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN30_N22190_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN30_N22190_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN30_N22190_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN32_N22192_io_in = {CBMux_IPIN32_N22192_io_in_hi,CBMux_IPIN32_N22192_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN32_N22192_io_config = configBlock_ioBundle_confOut[100:96]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN32_N22192_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN32_N22192_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN32_N22192_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN34_N22194_io_in = {CBMux_IPIN34_N22194_io_in_hi,CBMux_IPIN34_N22194_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN34_N22194_io_config = configBlock_ioBundle_confOut[105:101]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN34_N22194_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN34_N22194_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN34_N22194_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN36_N22196_io_in = {CBMux_IPIN36_N22196_io_in_hi,CBMux_IPIN36_N22196_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN36_N22196_io_config = configBlock_ioBundle_confOut[110:106]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN36_N22196_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN36_N22196_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN36_N22196_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN38_N22198_io_in = {CBMux_IPIN38_N22198_io_in_hi,CBMux_IPIN38_N22198_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN38_N22198_io_config = configBlock_ioBundle_confOut[115:111]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN38_N22198_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN38_N22198_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN38_N22198_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN40_N22200_io_in = {CBMux_IPIN40_N22200_io_in_hi,CBMux_IPIN40_N22200_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN40_N22200_io_config = configBlock_ioBundle_confOut[120:116]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN40_N22200_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN40_N22200_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN40_N22200_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN42_N22202_io_in = {CBMux_IPIN42_N22202_io_in_hi,CBMux_IPIN42_N22202_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN42_N22202_io_config = configBlock_ioBundle_confOut[125:121]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN42_N22202_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN42_N22202_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN42_N22202_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN44_N22204_io_in = {CBMux_IPIN44_N22204_io_in_hi,CBMux_IPIN44_N22204_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN44_N22204_io_config = configBlock_ioBundle_confOut[130:126]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN44_N22204_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN44_N22204_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN44_N22204_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN46_N22206_io_in = {CBMux_IPIN32_N22192_io_in_hi,CBMux_IPIN32_N22192_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN46_N22206_io_config = configBlock_ioBundle_confOut[135:131]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN46_N22206_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN46_N22206_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN46_N22206_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN48_N22208_io_in = {CBMux_IPIN40_N22200_io_in_hi,CBMux_IPIN40_N22200_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN48_N22208_io_config = configBlock_ioBundle_confOut[140:136]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN48_N22208_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN48_N22208_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN48_N22208_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN50_N22210_io_in = {CBMux_IPIN50_N22210_io_in_hi,CBMux_IPIN50_N22210_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN50_N22210_io_config = configBlock_ioBundle_confOut[145:141]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN50_N22210_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN50_N22210_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN50_N22210_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN52_N22212_io_in = {CBMux_IPIN36_N22196_io_in_hi,CBMux_IPIN36_N22196_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN52_N22212_io_config = configBlock_ioBundle_confOut[150:146]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN52_N22212_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN52_N22212_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN52_N22212_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN54_N22214_io_in = {CBMux_IPIN54_N22214_io_in_hi,CBMux_IPIN54_N22214_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN54_N22214_io_config = configBlock_ioBundle_confOut[155:151]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN54_N22214_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN54_N22214_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN54_N22214_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN56_N22216_io_in = {CBMux_IPIN56_N22216_io_in_hi,CBMux_IPIN56_N22216_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN56_N22216_io_config = configBlock_ioBundle_confOut[160:156]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN56_N22216_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN56_N22216_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN56_N22216_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN58_N22218_io_in = {CBMux_IPIN34_N22194_io_in_hi,CBMux_IPIN34_N22194_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN58_N22218_io_config = configBlock_ioBundle_confOut[165:161]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN58_N22218_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN58_N22218_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN58_N22218_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN60_N22220_io_in = {CBMux_IPIN42_N22202_io_in_hi,CBMux_IPIN42_N22202_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN60_N22220_io_config = configBlock_ioBundle_confOut[170:166]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN60_N22220_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN60_N22220_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN60_N22220_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN62_N22222_io_in = {CBMux_IPIN62_N22222_io_in_hi,CBMux_IPIN62_N22222_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN62_N22222_io_config = configBlock_ioBundle_confOut[175:171]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN62_N22222_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN62_N22222_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN62_N22222_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign SBMux_C5_N24197_O_7_C_1_io_in = {SBMux_C5_N24197_O_7_C_1_io_in_hi,SBMux_C5_N24197_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C5_N24197_O_7_C_1_io_config = configBlock_ioBundle_confOut[179:176]; // @[TileFull.scala 142:60]
  assign SBMux_C5_N24197_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C5_N24197_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C5_N24197_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C5_N24197_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C13_N24199_O_7_C_1_io_in = {SBMux_C13_N24199_O_7_C_1_io_in_hi,SBMux_C13_N24199_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C13_N24199_O_7_C_1_io_config = configBlock_ioBundle_confOut[183:180]; // @[TileFull.scala 142:60]
  assign SBMux_C13_N24199_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C13_N24199_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C13_N24199_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C13_N24199_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C21_N24201_O_7_C_1_io_in = {SBMux_C21_N24201_O_7_C_1_io_in_hi,SBMux_C21_N24201_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C21_N24201_O_7_C_1_io_config = configBlock_ioBundle_confOut[187:184]; // @[TileFull.scala 142:60]
  assign SBMux_C21_N24201_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C21_N24201_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C21_N24201_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C21_N24201_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C29_N24203_O_6_C_1_io_in = {SBMux_C29_N24203_O_6_C_1_io_in_hi,SBMux_C29_N24203_O_6_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C29_N24203_O_6_C_1_io_config = configBlock_ioBundle_confOut[191:188]; // @[TileFull.scala 142:60]
  assign SBMux_C29_N24203_O_6_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C29_N24203_O_6_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C29_N24203_O_6_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C29_N24203_O_6_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C37_N24205_O_6_C_2_io_in = {SBMux_C37_N24205_O_6_C_2_io_in_hi,SBMux_C37_N24205_O_6_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C37_N24205_O_6_C_2_io_config = configBlock_ioBundle_confOut[195:192]; // @[TileFull.scala 142:60]
  assign SBMux_C37_N24205_O_6_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C37_N24205_O_6_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C37_N24205_O_6_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C37_N24205_O_6_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C45_N24207_O_7_C_2_io_in = {SBMux_C45_N24207_O_7_C_2_io_in_hi,SBMux_C45_N24207_O_7_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C45_N24207_O_7_C_2_io_config = configBlock_ioBundle_confOut[199:196]; // @[TileFull.scala 142:60]
  assign SBMux_C45_N24207_O_7_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C45_N24207_O_7_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C45_N24207_O_7_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C45_N24207_O_7_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C53_N24209_O_7_C_1_io_in = {SBMux_C53_N24209_O_7_C_1_io_in_hi,SBMux_C53_N24209_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C53_N24209_O_7_C_1_io_config = configBlock_ioBundle_confOut[203:200]; // @[TileFull.scala 142:60]
  assign SBMux_C53_N24209_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C53_N24209_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C53_N24209_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C53_N24209_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C61_N24211_O_7_C_1_io_in = {SBMux_C61_N24211_O_7_C_1_io_in_hi,SBMux_C61_N24211_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C61_N24211_O_7_C_1_io_config = configBlock_ioBundle_confOut[207:204]; // @[TileFull.scala 142:60]
  assign SBMux_C61_N24211_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C61_N24211_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C61_N24211_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C61_N24211_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C69_N24213_O_6_C_1_io_in = {SBMux_C69_N24213_O_6_C_1_io_in_hi,SBMux_C29_N24203_O_6_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C69_N24213_O_6_C_1_io_config = configBlock_ioBundle_confOut[211:208]; // @[TileFull.scala 142:60]
  assign SBMux_C69_N24213_O_6_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C69_N24213_O_6_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C69_N24213_O_6_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C69_N24213_O_6_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C7_N24217_O_7_C_1_io_in = {SBMux_C7_N24217_O_7_C_1_io_in_hi,SBMux_C45_N24207_O_7_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C7_N24217_O_7_C_1_io_config = configBlock_ioBundle_confOut[215:212]; // @[TileFull.scala 142:60]
  assign SBMux_C7_N24217_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C7_N24217_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C7_N24217_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C7_N24217_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C15_N24219_O_7_C_1_io_in = {SBMux_C15_N24219_O_7_C_1_io_in_hi,SBMux_C53_N24209_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C15_N24219_O_7_C_1_io_config = configBlock_ioBundle_confOut[219:216]; // @[TileFull.scala 142:60]
  assign SBMux_C15_N24219_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C15_N24219_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C15_N24219_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C15_N24219_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C23_N24221_O_7_C_1_io_in = {SBMux_C23_N24221_O_7_C_1_io_in_hi,SBMux_C61_N24211_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C23_N24221_O_7_C_1_io_config = configBlock_ioBundle_confOut[223:220]; // @[TileFull.scala 142:60]
  assign SBMux_C23_N24221_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C23_N24221_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C23_N24221_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C23_N24221_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C31_N24223_O_6_C_1_io_in = {SBMux_C31_N24223_O_6_C_1_io_in_hi,SBMux_C29_N24203_O_6_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C31_N24223_O_6_C_1_io_config = configBlock_ioBundle_confOut[227:224]; // @[TileFull.scala 142:60]
  assign SBMux_C31_N24223_O_6_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C31_N24223_O_6_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C31_N24223_O_6_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C31_N24223_O_6_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C39_N24225_O_7_C_2_io_in = {SBMux_C39_N24225_O_7_C_2_io_in_hi,SBMux_C39_N24225_O_7_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C39_N24225_O_7_C_2_io_config = configBlock_ioBundle_confOut[231:228]; // @[TileFull.scala 142:60]
  assign SBMux_C39_N24225_O_7_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C39_N24225_O_7_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C39_N24225_O_7_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C39_N24225_O_7_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C47_N24227_O_7_C_2_io_in = {SBMux_C47_N24227_O_7_C_2_io_in_hi,SBMux_C47_N24227_O_7_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C47_N24227_O_7_C_2_io_config = configBlock_ioBundle_confOut[235:232]; // @[TileFull.scala 142:60]
  assign SBMux_C47_N24227_O_7_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C47_N24227_O_7_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C47_N24227_O_7_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C47_N24227_O_7_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C55_N24229_O_7_C_1_io_in = {SBMux_C55_N24229_O_7_C_1_io_in_hi,SBMux_C55_N24229_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C55_N24229_O_7_C_1_io_config = configBlock_ioBundle_confOut[239:236]; // @[TileFull.scala 142:60]
  assign SBMux_C55_N24229_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C55_N24229_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C55_N24229_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C55_N24229_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C63_N24231_O_7_C_1_io_in = {SBMux_C63_N24231_O_7_C_1_io_in_hi,SBMux_C63_N24231_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C63_N24231_O_7_C_1_io_config = configBlock_ioBundle_confOut[243:240]; // @[TileFull.scala 142:60]
  assign SBMux_C63_N24231_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C63_N24231_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C63_N24231_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C63_N24231_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C71_N24233_O_6_C_1_io_in = {SBMux_C71_N24233_O_6_C_1_io_in_hi,SBMux_C71_N24233_O_6_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C71_N24233_O_6_C_1_io_config = configBlock_ioBundle_confOut[247:244]; // @[TileFull.scala 142:60]
  assign SBMux_C71_N24233_O_6_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C71_N24233_O_6_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C71_N24233_O_6_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C71_N24233_O_6_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C1_N24237_O_7_C_1_io_in = {SBMux_C1_N24237_O_7_C_1_io_in_hi,SBMux_C39_N24225_O_7_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C1_N24237_O_7_C_1_io_config = configBlock_ioBundle_confOut[251:248]; // @[TileFull.scala 142:60]
  assign SBMux_C1_N24237_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C1_N24237_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C1_N24237_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C1_N24237_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C9_N24239_O_7_C_1_io_in = {SBMux_C9_N24239_O_7_C_1_io_in_hi,SBMux_C47_N24227_O_7_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C9_N24239_O_7_C_1_io_config = configBlock_ioBundle_confOut[255:252]; // @[TileFull.scala 142:60]
  assign SBMux_C9_N24239_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C9_N24239_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C9_N24239_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C9_N24239_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C17_N24241_O_7_C_1_io_in = {SBMux_C17_N24241_O_7_C_1_io_in_hi,SBMux_C55_N24229_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C17_N24241_O_7_C_1_io_config = configBlock_ioBundle_confOut[259:256]; // @[TileFull.scala 142:60]
  assign SBMux_C17_N24241_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C17_N24241_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C17_N24241_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C17_N24241_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C25_N24243_O_7_C_1_io_in = {SBMux_C25_N24243_O_7_C_1_io_in_hi,SBMux_C63_N24231_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C25_N24243_O_7_C_1_io_config = configBlock_ioBundle_confOut[263:260]; // @[TileFull.scala 142:60]
  assign SBMux_C25_N24243_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C25_N24243_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C25_N24243_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C25_N24243_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C33_N24245_O_6_C_1_io_in = {SBMux_C33_N24245_O_6_C_1_io_in_hi,SBMux_C71_N24233_O_6_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C33_N24245_O_6_C_1_io_config = configBlock_ioBundle_confOut[267:264]; // @[TileFull.scala 142:60]
  assign SBMux_C33_N24245_O_6_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C33_N24245_O_6_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C33_N24245_O_6_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C33_N24245_O_6_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C41_N24247_O_7_C_2_io_in = {SBMux_C41_N24247_O_7_C_2_io_in_hi,SBMux_C41_N24247_O_7_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C41_N24247_O_7_C_2_io_config = configBlock_ioBundle_confOut[271:268]; // @[TileFull.scala 142:60]
  assign SBMux_C41_N24247_O_7_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C41_N24247_O_7_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C41_N24247_O_7_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C41_N24247_O_7_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C49_N24249_O_7_C_2_io_in = {SBMux_C49_N24249_O_7_C_2_io_in_hi,SBMux_C49_N24249_O_7_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C49_N24249_O_7_C_2_io_config = configBlock_ioBundle_confOut[275:272]; // @[TileFull.scala 142:60]
  assign SBMux_C49_N24249_O_7_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C49_N24249_O_7_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C49_N24249_O_7_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C49_N24249_O_7_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C57_N24251_O_7_C_1_io_in = {SBMux_C57_N24251_O_7_C_1_io_in_hi,SBMux_C57_N24251_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C57_N24251_O_7_C_1_io_config = configBlock_ioBundle_confOut[279:276]; // @[TileFull.scala 142:60]
  assign SBMux_C57_N24251_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C57_N24251_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C57_N24251_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C57_N24251_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C65_N24253_O_7_C_1_io_in = {SBMux_C65_N24253_O_7_C_1_io_in_hi,SBMux_C65_N24253_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C65_N24253_O_7_C_1_io_config = configBlock_ioBundle_confOut[283:280]; // @[TileFull.scala 142:60]
  assign SBMux_C65_N24253_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C65_N24253_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C65_N24253_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C65_N24253_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C73_N24255_O_6_C_1_io_in = {SBMux_C73_N24255_O_6_C_1_io_in_hi,SBMux_C73_N24255_O_6_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C73_N24255_O_6_C_1_io_config = configBlock_ioBundle_confOut[287:284]; // @[TileFull.scala 142:60]
  assign SBMux_C73_N24255_O_6_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C73_N24255_O_6_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C73_N24255_O_6_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C73_N24255_O_6_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C77_N24257_O_16_C_1_io_in = {SBMux_C77_N24257_O_16_C_1_io_in_hi,SBMux_C77_N24257_O_16_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C77_N24257_O_16_C_1_io_config = configBlock_ioBundle_confOut[292:288]; // @[TileFull.scala 142:60]
  assign SBMux_C77_N24257_O_16_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C77_N24257_O_16_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C77_N24257_O_16_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C77_N24257_O_16_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C3_N24259_O_7_C_1_io_in = {SBMux_C3_N24259_O_7_C_1_io_in_hi,SBMux_C41_N24247_O_7_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C3_N24259_O_7_C_1_io_config = configBlock_ioBundle_confOut[296:293]; // @[TileFull.scala 142:60]
  assign SBMux_C3_N24259_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C3_N24259_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C3_N24259_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C3_N24259_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C11_N24261_O_7_C_1_io_in = {SBMux_C11_N24261_O_7_C_1_io_in_hi,SBMux_C49_N24249_O_7_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C11_N24261_O_7_C_1_io_config = configBlock_ioBundle_confOut[300:297]; // @[TileFull.scala 142:60]
  assign SBMux_C11_N24261_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C11_N24261_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C11_N24261_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C11_N24261_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C19_N24263_O_7_C_1_io_in = {SBMux_C19_N24263_O_7_C_1_io_in_hi,SBMux_C57_N24251_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C19_N24263_O_7_C_1_io_config = configBlock_ioBundle_confOut[304:301]; // @[TileFull.scala 142:60]
  assign SBMux_C19_N24263_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C19_N24263_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C19_N24263_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C19_N24263_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C27_N24265_O_7_C_1_io_in = {SBMux_C27_N24265_O_7_C_1_io_in_hi,SBMux_C65_N24253_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C27_N24265_O_7_C_1_io_config = configBlock_ioBundle_confOut[308:305]; // @[TileFull.scala 142:60]
  assign SBMux_C27_N24265_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C27_N24265_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C27_N24265_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C27_N24265_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C35_N24267_O_6_C_2_io_in = {SBMux_C35_N24267_O_6_C_2_io_in_hi,SBMux_C35_N24267_O_6_C_2_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C35_N24267_O_6_C_2_io_config = configBlock_ioBundle_confOut[312:309]; // @[TileFull.scala 142:60]
  assign SBMux_C35_N24267_O_6_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C35_N24267_O_6_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C35_N24267_O_6_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C35_N24267_O_6_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C43_N24269_O_7_C_2_io_in = {SBMux_C43_N24269_O_7_C_2_io_in_hi,SBMux_C5_N24197_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C43_N24269_O_7_C_2_io_config = configBlock_ioBundle_confOut[316:313]; // @[TileFull.scala 142:60]
  assign SBMux_C43_N24269_O_7_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C43_N24269_O_7_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C43_N24269_O_7_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C43_N24269_O_7_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C51_N24271_O_7_C_1_io_in = {SBMux_C51_N24271_O_7_C_1_io_in_hi,SBMux_C13_N24199_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C51_N24271_O_7_C_1_io_config = configBlock_ioBundle_confOut[320:317]; // @[TileFull.scala 142:60]
  assign SBMux_C51_N24271_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C51_N24271_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C51_N24271_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C51_N24271_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C59_N24273_O_7_C_1_io_in = {SBMux_C59_N24273_O_7_C_1_io_in_hi,SBMux_C21_N24201_O_7_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C59_N24273_O_7_C_1_io_config = configBlock_ioBundle_confOut[324:321]; // @[TileFull.scala 142:60]
  assign SBMux_C59_N24273_O_7_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C59_N24273_O_7_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C59_N24273_O_7_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C59_N24273_O_7_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C67_N24275_O_6_C_1_io_in = {SBMux_C67_N24275_O_6_C_1_io_in_hi,SBMux_C29_N24203_O_6_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C67_N24275_O_6_C_1_io_config = configBlock_ioBundle_confOut[328:325]; // @[TileFull.scala 142:60]
  assign SBMux_C67_N24275_O_6_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C67_N24275_O_6_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C67_N24275_O_6_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C67_N24275_O_6_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C75_N24277_O_6_C_1_io_in = {SBMux_C75_N24277_O_6_C_1_io_in_hi,SBMux_C75_N24277_O_6_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C75_N24277_O_6_C_1_io_config = configBlock_ioBundle_confOut[332:329]; // @[TileFull.scala 142:60]
  assign SBMux_C75_N24277_O_6_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C75_N24277_O_6_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C75_N24277_O_6_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C75_N24277_O_6_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C79_N24279_O_16_C_1_io_in = {SBMux_C79_N24279_O_16_C_1_io_in_hi,SBMux_C79_N24279_O_16_C_1_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C79_N24279_O_16_C_1_io_config = configBlock_ioBundle_confOut[337:333]; // @[TileFull.scala 142:60]
  assign SBMux_C79_N24279_O_16_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C79_N24279_O_16_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C79_N24279_O_16_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C79_N24279_O_16_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C5_N29271_O_0_C_5_io_in = {SBMux_C5_N29271_O_0_C_5_io_in_hi,SBMux_C5_N29271_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C5_N29271_O_0_C_5_io_config = configBlock_ioBundle_confOut[341:338]; // @[TileFull.scala 142:60]
  assign SBMux_C5_N29271_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C5_N29271_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C5_N29271_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C5_N29271_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C13_N29279_O_0_C_5_io_in = {SBMux_C13_N29279_O_0_C_5_io_in_hi,SBMux_C13_N29279_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C13_N29279_O_0_C_5_io_config = configBlock_ioBundle_confOut[345:342]; // @[TileFull.scala 142:60]
  assign SBMux_C13_N29279_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C13_N29279_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C13_N29279_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C13_N29279_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C21_N29287_O_0_C_5_io_in = {SBMux_C21_N29287_O_0_C_5_io_in_hi,SBMux_C21_N29287_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C21_N29287_O_0_C_5_io_config = configBlock_ioBundle_confOut[349:346]; // @[TileFull.scala 142:60]
  assign SBMux_C21_N29287_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C21_N29287_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C21_N29287_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C21_N29287_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C29_N29295_O_0_C_5_io_in = {SBMux_C29_N29295_O_0_C_5_io_in_hi,SBMux_C29_N29295_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C29_N29295_O_0_C_5_io_config = configBlock_ioBundle_confOut[353:350]; // @[TileFull.scala 142:60]
  assign SBMux_C29_N29295_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C29_N29295_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C29_N29295_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C29_N29295_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C37_N29303_O_0_C_5_io_in = {SBMux_C37_N29303_O_0_C_5_io_in_hi,SBMux_C37_N29303_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C37_N29303_O_0_C_5_io_config = configBlock_ioBundle_confOut[357:354]; // @[TileFull.scala 142:60]
  assign SBMux_C37_N29303_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C37_N29303_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C37_N29303_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C37_N29303_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C45_N29311_O_0_C_5_io_in = {SBMux_C45_N29311_O_0_C_5_io_in_hi,SBMux_C45_N29311_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C45_N29311_O_0_C_5_io_config = configBlock_ioBundle_confOut[361:358]; // @[TileFull.scala 142:60]
  assign SBMux_C45_N29311_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C45_N29311_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C45_N29311_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C45_N29311_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C53_N29319_O_0_C_5_io_in = {SBMux_C53_N29319_O_0_C_5_io_in_hi,SBMux_C53_N29319_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C53_N29319_O_0_C_5_io_config = configBlock_ioBundle_confOut[365:362]; // @[TileFull.scala 142:60]
  assign SBMux_C53_N29319_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C53_N29319_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C53_N29319_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C53_N29319_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C61_N29327_O_0_C_5_io_in = {SBMux_C61_N29327_O_0_C_5_io_in_hi,SBMux_C61_N29327_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C61_N29327_O_0_C_5_io_config = configBlock_ioBundle_confOut[369:366]; // @[TileFull.scala 142:60]
  assign SBMux_C61_N29327_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C61_N29327_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C61_N29327_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C61_N29327_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C69_N29335_O_0_C_5_io_in = {SBMux_C69_N29335_O_0_C_5_io_in_hi,SBMux_C69_N29335_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C69_N29335_O_0_C_5_io_config = configBlock_ioBundle_confOut[373:370]; // @[TileFull.scala 142:60]
  assign SBMux_C69_N29335_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C69_N29335_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C69_N29335_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C69_N29335_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C77_N29367_O_0_C_5_io_in = {SBMux_C77_N29367_O_0_C_5_io_in_hi,SBMux_C77_N29367_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C77_N29367_O_0_C_5_io_config = configBlock_ioBundle_confOut[377:374]; // @[TileFull.scala 142:60]
  assign SBMux_C77_N29367_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C77_N29367_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C77_N29367_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C77_N29367_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C4_N29390_O_0_C_5_io_in = {SBMux_C4_N29390_O_0_C_5_io_in_hi,SBMux_C77_N29367_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C4_N29390_O_0_C_5_io_config = configBlock_ioBundle_confOut[381:378]; // @[TileFull.scala 142:60]
  assign SBMux_C4_N29390_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C4_N29390_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C4_N29390_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C4_N29390_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C12_N29392_O_0_C_5_io_in = {SBMux_C12_N29392_O_0_C_5_io_in_hi,SBMux_C69_N29335_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C12_N29392_O_0_C_5_io_config = configBlock_ioBundle_confOut[385:382]; // @[TileFull.scala 142:60]
  assign SBMux_C12_N29392_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C12_N29392_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C12_N29392_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C12_N29392_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C20_N29394_O_0_C_5_io_in = {SBMux_C20_N29394_O_0_C_5_io_in_hi,SBMux_C61_N29327_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C20_N29394_O_0_C_5_io_config = configBlock_ioBundle_confOut[389:386]; // @[TileFull.scala 142:60]
  assign SBMux_C20_N29394_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C20_N29394_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C20_N29394_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C20_N29394_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C28_N29396_O_0_C_5_io_in = {SBMux_C28_N29396_O_0_C_5_io_in_hi,SBMux_C53_N29319_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C28_N29396_O_0_C_5_io_config = configBlock_ioBundle_confOut[393:390]; // @[TileFull.scala 142:60]
  assign SBMux_C28_N29396_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C28_N29396_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C28_N29396_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C28_N29396_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C36_N29398_O_0_C_5_io_in = {SBMux_C36_N29398_O_0_C_5_io_in_hi,SBMux_C45_N29311_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C36_N29398_O_0_C_5_io_config = configBlock_ioBundle_confOut[397:394]; // @[TileFull.scala 142:60]
  assign SBMux_C36_N29398_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C36_N29398_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C36_N29398_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C36_N29398_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C44_N29400_O_0_C_5_io_in = {SBMux_C44_N29400_O_0_C_5_io_in_hi,SBMux_C37_N29303_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C44_N29400_O_0_C_5_io_config = configBlock_ioBundle_confOut[401:398]; // @[TileFull.scala 142:60]
  assign SBMux_C44_N29400_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C44_N29400_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C44_N29400_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C44_N29400_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C52_N29402_O_0_C_5_io_in = {SBMux_C52_N29402_O_0_C_5_io_in_hi,SBMux_C29_N29295_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C52_N29402_O_0_C_5_io_config = configBlock_ioBundle_confOut[405:402]; // @[TileFull.scala 142:60]
  assign SBMux_C52_N29402_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C52_N29402_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C52_N29402_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C52_N29402_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C60_N29404_O_0_C_5_io_in = {SBMux_C60_N29404_O_0_C_5_io_in_hi,SBMux_C21_N29287_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C60_N29404_O_0_C_5_io_config = configBlock_ioBundle_confOut[409:406]; // @[TileFull.scala 142:60]
  assign SBMux_C60_N29404_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C60_N29404_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C60_N29404_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C60_N29404_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C68_N29406_O_0_C_5_io_in = {SBMux_C68_N29406_O_0_C_5_io_in_hi,SBMux_C13_N29279_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C68_N29406_O_0_C_5_io_config = configBlock_ioBundle_confOut[413:410]; // @[TileFull.scala 142:60]
  assign SBMux_C68_N29406_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C68_N29406_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C68_N29406_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C68_N29406_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C76_N29408_O_0_C_5_io_in = {SBMux_C76_N29408_O_0_C_5_io_in_hi,SBMux_C5_N29271_O_0_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C76_N29408_O_0_C_5_io_config = configBlock_ioBundle_confOut[417:414]; // @[TileFull.scala 142:60]
  assign SBMux_C76_N29408_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C76_N29408_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C76_N29408_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C76_N29408_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
endmodule
