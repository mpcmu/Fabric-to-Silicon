module Ble4(
  input         clock,
  input         reset,
  input  [19:0] io_config,
  input         io_in_0,
  input         io_in_1,
  input         io_in_2,
  input         io_in_3,
  output        io_outR,
  output        io_outT,
  input         io_gndOuts,
  input         io_clkEnb
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] lut_in; // @[CLBlut4N10Clb.scala 73:27]
  wire [3:0] lut_sel; // @[CLBlut4N10Clb.scala 73:27]
  wire  lut_o; // @[CLBlut4N10Clb.scala 73:27]
  wire [1:0] lut_io_sel_lo = {io_in_1,io_in_0}; // @[CLBlut4N10Clb.scala 75:23]
  wire [1:0] lut_io_sel_hi = {io_in_3,io_in_2}; // @[CLBlut4N10Clb.scala 75:23]
  wire  _bleFF_T = ~io_clkEnb; // @[CLBlut4N10Clb.scala 77:48]
  reg  bleFF; // @[Reg.scala 28:20]
  wire  _io_outR_T_1 = io_config[16] ? lut_o : bleFF; // @[CLBlut4N10Clb.scala 80:17]
  wire  _io_outR_T_2 = ~io_gndOuts; // @[CLBlut4N10Clb.scala 80:52]
  wire  _io_outT_T_1 = io_config[17] ? lut_o : bleFF; // @[CLBlut4N10Clb.scala 81:17]
  Mux16C lut ( // @[CLBlut4N10Clb.scala 73:27]
    .in(lut_in),
    .sel(lut_sel),
    .o(lut_o)
  );
  assign io_outR = _io_outR_T_1 & ~io_gndOuts; // @[CLBlut4N10Clb.scala 80:50]
  assign io_outT = _io_outT_T_1 & _io_outR_T_2; // @[CLBlut4N10Clb.scala 81:50]
  assign lut_in = io_config[15:0]; // @[CLBlut4N10Clb.scala 74:25]
  assign lut_sel = {lut_io_sel_hi,lut_io_sel_lo}; // @[CLBlut4N10Clb.scala 75:23]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      bleFF <= 1'h0; // @[Reg.scala 28:20]
    end else if (_bleFF_T) begin // @[Reg.scala 29:18]
      bleFF <= lut_o; // @[Reg.scala 29:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bleFF = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLBlut4N10Mem(
  input          IPIN_0,
  input          IPIN_1,
  input          IPIN_2,
  input          IPIN_3,
  input          IPIN_4,
  input          IPIN_5,
  input          IPIN_6,
  input          IPIN_7,
  input          IPIN_8,
  input          IPIN_9,
  input          IPIN_10,
  input          IPIN_11,
  input          IPIN_12,
  input          IPIN_13,
  input          IPIN_14,
  input          IPIN_15,
  input          IPIN_16,
  input          IPIN_17,
  input          IPIN_18,
  input          IPIN_19,
  input          IPIN_20,
  input          IPIN_21,
  input          IPIN_22,
  input          IPIN_23,
  input          IPIN_24,
  input          IPIN_25,
  input          IPIN_26,
  input          IPIN_27,
  input          IPIN_28,
  input          IPIN_29,
  input          IPIN_30,
  input          IPIN_31,
  output         OPIN_41,
  output         OPIN_42,
  output         OPIN_43,
  output         OPIN_44,
  output         OPIN_45,
  output         OPIN_46,
  output         OPIN_47,
  output         OPIN_48,
  output         OPIN_49,
  output         OPIN_50,
  output         OPIN_51,
  output         OPIN_52,
  output         OPIN_53,
  output         OPIN_54,
  output         OPIN_55,
  output         OPIN_56,
  input          clock,
  input          reset,
  input  [15:0]  ioPad_i,
  input  [161:0] configBits,
  input          gndLBouts
);
  wire  BLE_0_clock; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_0_reset; // @[CLBlut4N10Mem.scala 54:48]
  wire [19:0] BLE_0_io_config; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_0_io_in_0; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_0_io_in_1; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_0_io_in_2; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_0_io_in_3; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_0_io_outR; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_0_io_outT; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_0_io_gndOuts; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_0_io_clkEnb; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_1_clock; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_1_reset; // @[CLBlut4N10Mem.scala 54:48]
  wire [19:0] BLE_1_io_config; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_1_io_in_0; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_1_io_in_1; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_1_io_in_2; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_1_io_in_3; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_1_io_outR; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_1_io_outT; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_1_io_gndOuts; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_1_io_clkEnb; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_2_clock; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_2_reset; // @[CLBlut4N10Mem.scala 54:48]
  wire [19:0] BLE_2_io_config; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_2_io_in_0; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_2_io_in_1; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_2_io_in_2; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_2_io_in_3; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_2_io_outR; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_2_io_outT; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_2_io_gndOuts; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_2_io_clkEnb; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_3_clock; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_3_reset; // @[CLBlut4N10Mem.scala 54:48]
  wire [19:0] BLE_3_io_config; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_3_io_in_0; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_3_io_in_1; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_3_io_in_2; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_3_io_in_3; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_3_io_outR; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_3_io_outT; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_3_io_gndOuts; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_3_io_clkEnb; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_4_clock; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_4_reset; // @[CLBlut4N10Mem.scala 54:48]
  wire [19:0] BLE_4_io_config; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_4_io_in_0; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_4_io_in_1; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_4_io_in_2; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_4_io_in_3; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_4_io_outR; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_4_io_outT; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_4_io_gndOuts; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_4_io_clkEnb; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_5_clock; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_5_reset; // @[CLBlut4N10Mem.scala 54:48]
  wire [19:0] BLE_5_io_config; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_5_io_in_0; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_5_io_in_1; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_5_io_in_2; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_5_io_in_3; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_5_io_outR; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_5_io_outT; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_5_io_gndOuts; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_5_io_clkEnb; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_6_clock; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_6_reset; // @[CLBlut4N10Mem.scala 54:48]
  wire [19:0] BLE_6_io_config; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_6_io_in_0; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_6_io_in_1; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_6_io_in_2; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_6_io_in_3; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_6_io_outR; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_6_io_outT; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_6_io_gndOuts; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_6_io_clkEnb; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_7_clock; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_7_reset; // @[CLBlut4N10Mem.scala 54:48]
  wire [19:0] BLE_7_io_config; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_7_io_in_0; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_7_io_in_1; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_7_io_in_2; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_7_io_in_3; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_7_io_outR; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_7_io_outT; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_7_io_gndOuts; // @[CLBlut4N10Mem.scala 54:48]
  wire  BLE_7_io_clkEnb; // @[CLBlut4N10Mem.scala 54:48]
  wire [7:0] I_0 = {IPIN_7,IPIN_6,IPIN_5,IPIN_4,IPIN_3,IPIN_2,IPIN_1,IPIN_0}; // @[CLBlut4N10Mem.scala 35:92]
  wire [7:0] I_1 = {IPIN_15,IPIN_14,IPIN_13,IPIN_12,IPIN_11,IPIN_10,IPIN_9,IPIN_8}; // @[CLBlut4N10Mem.scala 35:92]
  wire [7:0] I_2 = {IPIN_23,IPIN_22,IPIN_21,IPIN_20,IPIN_19,IPIN_18,IPIN_17,IPIN_16}; // @[CLBlut4N10Mem.scala 35:92]
  wire [7:0] I_3 = {IPIN_31,IPIN_30,IPIN_29,IPIN_28,IPIN_27,IPIN_26,IPIN_25,IPIN_24}; // @[CLBlut4N10Mem.scala 35:92]
  wire  OMem_0 = ioPad_i[0]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_0 = BLE_0_io_outR; // @[CLBlut4N10Mem.scala 38:18 58:15]
  wire  OMem_1 = ioPad_i[1]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_1 = BLE_1_io_outR; // @[CLBlut4N10Mem.scala 38:18 58:15]
  wire  OMem_2 = ioPad_i[2]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_2 = BLE_2_io_outR; // @[CLBlut4N10Mem.scala 38:18 58:15]
  wire  OMem_3 = ioPad_i[3]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_3 = BLE_3_io_outR; // @[CLBlut4N10Mem.scala 38:18 58:15]
  wire  OMem_4 = ioPad_i[4]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_4 = BLE_4_io_outR; // @[CLBlut4N10Mem.scala 38:18 58:15]
  wire  OMem_5 = ioPad_i[5]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_5 = BLE_5_io_outR; // @[CLBlut4N10Mem.scala 38:18 58:15]
  wire  OMem_6 = ioPad_i[6]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_6 = BLE_6_io_outR; // @[CLBlut4N10Mem.scala 38:18 58:15]
  wire  OMem_7 = ioPad_i[7]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_7 = BLE_7_io_outR; // @[CLBlut4N10Mem.scala 38:18 58:15]
  wire  OMem_8 = ioPad_i[8]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_8 = BLE_0_io_outT; // @[CLBlut4N10Mem.scala 38:18 59:17]
  wire  OMem_9 = ioPad_i[9]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_9 = BLE_1_io_outT; // @[CLBlut4N10Mem.scala 38:18 59:17]
  wire  OMem_10 = ioPad_i[10]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_10 = BLE_2_io_outT; // @[CLBlut4N10Mem.scala 38:18 59:17]
  wire  OMem_11 = ioPad_i[11]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_11 = BLE_3_io_outT; // @[CLBlut4N10Mem.scala 38:18 59:17]
  wire  OMem_12 = ioPad_i[12]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_12 = BLE_4_io_outT; // @[CLBlut4N10Mem.scala 38:18 59:17]
  wire  OMem_13 = ioPad_i[13]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_13 = BLE_5_io_outT; // @[CLBlut4N10Mem.scala 38:18 59:17]
  wire  OMem_14 = ioPad_i[14]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_14 = BLE_6_io_outT; // @[CLBlut4N10Mem.scala 38:18 59:17]
  wire  OMem_15 = ioPad_i[15]; // @[CLBlut4N10Mem.scala 47:65]
  wire  OClb_15 = BLE_7_io_outT; // @[CLBlut4N10Mem.scala 38:18 59:17]
  Ble4 BLE_0 ( // @[CLBlut4N10Mem.scala 54:48]
    .clock(BLE_0_clock),
    .reset(BLE_0_reset),
    .io_config(BLE_0_io_config),
    .io_in_0(BLE_0_io_in_0),
    .io_in_1(BLE_0_io_in_1),
    .io_in_2(BLE_0_io_in_2),
    .io_in_3(BLE_0_io_in_3),
    .io_outR(BLE_0_io_outR),
    .io_outT(BLE_0_io_outT),
    .io_gndOuts(BLE_0_io_gndOuts),
    .io_clkEnb(BLE_0_io_clkEnb)
  );
  Ble4 BLE_1 ( // @[CLBlut4N10Mem.scala 54:48]
    .clock(BLE_1_clock),
    .reset(BLE_1_reset),
    .io_config(BLE_1_io_config),
    .io_in_0(BLE_1_io_in_0),
    .io_in_1(BLE_1_io_in_1),
    .io_in_2(BLE_1_io_in_2),
    .io_in_3(BLE_1_io_in_3),
    .io_outR(BLE_1_io_outR),
    .io_outT(BLE_1_io_outT),
    .io_gndOuts(BLE_1_io_gndOuts),
    .io_clkEnb(BLE_1_io_clkEnb)
  );
  Ble4 BLE_2 ( // @[CLBlut4N10Mem.scala 54:48]
    .clock(BLE_2_clock),
    .reset(BLE_2_reset),
    .io_config(BLE_2_io_config),
    .io_in_0(BLE_2_io_in_0),
    .io_in_1(BLE_2_io_in_1),
    .io_in_2(BLE_2_io_in_2),
    .io_in_3(BLE_2_io_in_3),
    .io_outR(BLE_2_io_outR),
    .io_outT(BLE_2_io_outT),
    .io_gndOuts(BLE_2_io_gndOuts),
    .io_clkEnb(BLE_2_io_clkEnb)
  );
  Ble4 BLE_3 ( // @[CLBlut4N10Mem.scala 54:48]
    .clock(BLE_3_clock),
    .reset(BLE_3_reset),
    .io_config(BLE_3_io_config),
    .io_in_0(BLE_3_io_in_0),
    .io_in_1(BLE_3_io_in_1),
    .io_in_2(BLE_3_io_in_2),
    .io_in_3(BLE_3_io_in_3),
    .io_outR(BLE_3_io_outR),
    .io_outT(BLE_3_io_outT),
    .io_gndOuts(BLE_3_io_gndOuts),
    .io_clkEnb(BLE_3_io_clkEnb)
  );
  Ble4 BLE_4 ( // @[CLBlut4N10Mem.scala 54:48]
    .clock(BLE_4_clock),
    .reset(BLE_4_reset),
    .io_config(BLE_4_io_config),
    .io_in_0(BLE_4_io_in_0),
    .io_in_1(BLE_4_io_in_1),
    .io_in_2(BLE_4_io_in_2),
    .io_in_3(BLE_4_io_in_3),
    .io_outR(BLE_4_io_outR),
    .io_outT(BLE_4_io_outT),
    .io_gndOuts(BLE_4_io_gndOuts),
    .io_clkEnb(BLE_4_io_clkEnb)
  );
  Ble4 BLE_5 ( // @[CLBlut4N10Mem.scala 54:48]
    .clock(BLE_5_clock),
    .reset(BLE_5_reset),
    .io_config(BLE_5_io_config),
    .io_in_0(BLE_5_io_in_0),
    .io_in_1(BLE_5_io_in_1),
    .io_in_2(BLE_5_io_in_2),
    .io_in_3(BLE_5_io_in_3),
    .io_outR(BLE_5_io_outR),
    .io_outT(BLE_5_io_outT),
    .io_gndOuts(BLE_5_io_gndOuts),
    .io_clkEnb(BLE_5_io_clkEnb)
  );
  Ble4 BLE_6 ( // @[CLBlut4N10Mem.scala 54:48]
    .clock(BLE_6_clock),
    .reset(BLE_6_reset),
    .io_config(BLE_6_io_config),
    .io_in_0(BLE_6_io_in_0),
    .io_in_1(BLE_6_io_in_1),
    .io_in_2(BLE_6_io_in_2),
    .io_in_3(BLE_6_io_in_3),
    .io_outR(BLE_6_io_outR),
    .io_outT(BLE_6_io_outT),
    .io_gndOuts(BLE_6_io_gndOuts),
    .io_clkEnb(BLE_6_io_clkEnb)
  );
  Ble4 BLE_7 ( // @[CLBlut4N10Mem.scala 54:48]
    .clock(BLE_7_clock),
    .reset(BLE_7_reset),
    .io_config(BLE_7_io_config),
    .io_in_0(BLE_7_io_in_0),
    .io_in_1(BLE_7_io_in_1),
    .io_in_2(BLE_7_io_in_2),
    .io_in_3(BLE_7_io_in_3),
    .io_outR(BLE_7_io_outR),
    .io_outT(BLE_7_io_outT),
    .io_gndOuts(BLE_7_io_gndOuts),
    .io_clkEnb(BLE_7_io_clkEnb)
  );
  assign OPIN_41 = configBits[160] ? OMem_0 : OClb_0; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_42 = configBits[160] ? OMem_1 : OClb_1; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_43 = configBits[160] ? OMem_2 : OClb_2; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_44 = configBits[160] ? OMem_3 : OClb_3; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_45 = configBits[160] ? OMem_4 : OClb_4; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_46 = configBits[160] ? OMem_5 : OClb_5; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_47 = configBits[160] ? OMem_6 : OClb_6; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_48 = configBits[160] ? OMem_7 : OClb_7; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_49 = configBits[160] ? OMem_8 : OClb_8; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_50 = configBits[160] ? OMem_9 : OClb_9; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_51 = configBits[160] ? OMem_10 : OClb_10; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_52 = configBits[160] ? OMem_11 : OClb_11; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_53 = configBits[160] ? OMem_12 : OClb_12; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_54 = configBits[160] ? OMem_13 : OClb_13; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_55 = configBits[160] ? OMem_14 : OClb_14; // @[CLBlut4N10Mem.scala 40:15]
  assign OPIN_56 = configBits[160] ? OMem_15 : OClb_15; // @[CLBlut4N10Mem.scala 40:15]
  assign BLE_0_clock = clock;
  assign BLE_0_reset = reset;
  assign BLE_0_io_config = configBits[19:0]; // @[CLBlut4N10Mem.scala 56:38]
  assign BLE_0_io_in_0 = I_0[0]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_0_io_in_1 = I_1[0]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_0_io_in_2 = I_2[0]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_0_io_in_3 = I_3[0]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_0_io_gndOuts = gndLBouts; // @[CLBlut4N10Mem.scala 60:26]
  assign BLE_0_io_clkEnb = configBits[161]; // @[CLBlut4N10Mem.scala 61:38]
  assign BLE_1_clock = clock;
  assign BLE_1_reset = reset;
  assign BLE_1_io_config = configBits[39:20]; // @[CLBlut4N10Mem.scala 56:38]
  assign BLE_1_io_in_0 = I_0[1]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_1_io_in_1 = I_1[1]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_1_io_in_2 = I_2[1]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_1_io_in_3 = I_3[1]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_1_io_gndOuts = gndLBouts; // @[CLBlut4N10Mem.scala 60:26]
  assign BLE_1_io_clkEnb = configBits[161]; // @[CLBlut4N10Mem.scala 61:38]
  assign BLE_2_clock = clock;
  assign BLE_2_reset = reset;
  assign BLE_2_io_config = configBits[59:40]; // @[CLBlut4N10Mem.scala 56:38]
  assign BLE_2_io_in_0 = I_0[2]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_2_io_in_1 = I_1[2]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_2_io_in_2 = I_2[2]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_2_io_in_3 = I_3[2]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_2_io_gndOuts = gndLBouts; // @[CLBlut4N10Mem.scala 60:26]
  assign BLE_2_io_clkEnb = configBits[161]; // @[CLBlut4N10Mem.scala 61:38]
  assign BLE_3_clock = clock;
  assign BLE_3_reset = reset;
  assign BLE_3_io_config = configBits[79:60]; // @[CLBlut4N10Mem.scala 56:38]
  assign BLE_3_io_in_0 = I_0[3]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_3_io_in_1 = I_1[3]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_3_io_in_2 = I_2[3]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_3_io_in_3 = I_3[3]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_3_io_gndOuts = gndLBouts; // @[CLBlut4N10Mem.scala 60:26]
  assign BLE_3_io_clkEnb = configBits[161]; // @[CLBlut4N10Mem.scala 61:38]
  assign BLE_4_clock = clock;
  assign BLE_4_reset = reset;
  assign BLE_4_io_config = configBits[99:80]; // @[CLBlut4N10Mem.scala 56:38]
  assign BLE_4_io_in_0 = I_0[4]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_4_io_in_1 = I_1[4]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_4_io_in_2 = I_2[4]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_4_io_in_3 = I_3[4]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_4_io_gndOuts = gndLBouts; // @[CLBlut4N10Mem.scala 60:26]
  assign BLE_4_io_clkEnb = configBits[161]; // @[CLBlut4N10Mem.scala 61:38]
  assign BLE_5_clock = clock;
  assign BLE_5_reset = reset;
  assign BLE_5_io_config = configBits[119:100]; // @[CLBlut4N10Mem.scala 56:38]
  assign BLE_5_io_in_0 = I_0[5]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_5_io_in_1 = I_1[5]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_5_io_in_2 = I_2[5]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_5_io_in_3 = I_3[5]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_5_io_gndOuts = gndLBouts; // @[CLBlut4N10Mem.scala 60:26]
  assign BLE_5_io_clkEnb = configBits[161]; // @[CLBlut4N10Mem.scala 61:38]
  assign BLE_6_clock = clock;
  assign BLE_6_reset = reset;
  assign BLE_6_io_config = configBits[139:120]; // @[CLBlut4N10Mem.scala 56:38]
  assign BLE_6_io_in_0 = I_0[6]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_6_io_in_1 = I_1[6]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_6_io_in_2 = I_2[6]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_6_io_in_3 = I_3[6]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_6_io_gndOuts = gndLBouts; // @[CLBlut4N10Mem.scala 60:26]
  assign BLE_6_io_clkEnb = configBits[161]; // @[CLBlut4N10Mem.scala 61:38]
  assign BLE_7_clock = clock;
  assign BLE_7_reset = reset;
  assign BLE_7_io_config = configBits[159:140]; // @[CLBlut4N10Mem.scala 56:38]
  assign BLE_7_io_in_0 = I_0[7]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_7_io_in_1 = I_1[7]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_7_io_in_2 = I_2[7]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_7_io_in_3 = I_3[7]; // @[CLBlut4N10Mem.scala 57:62]
  assign BLE_7_io_gndOuts = gndLBouts; // @[CLBlut4N10Mem.scala 60:26]
  assign BLE_7_io_clkEnb = configBits[161]; // @[CLBlut4N10Mem.scala 61:38]
endmodule
module ScanConf_Tile_9_3_clbmemtile(
  input          clock,
  output [495:0] ioBundle_confOut,
  input  [7:0]   ioBundle_scan_in,
  input          ioBundle_scan_en,
  output [7:0]   ioBundle_scan_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
`endif // RANDOMIZE_REG_INIT
  reg  confReg_0; // @[ScanConf.scala 32:20]
  reg  confReg_1; // @[ScanConf.scala 32:20]
  reg  confReg_2; // @[ScanConf.scala 32:20]
  reg  confReg_3; // @[ScanConf.scala 32:20]
  reg  confReg_4; // @[ScanConf.scala 32:20]
  reg  confReg_5; // @[ScanConf.scala 32:20]
  reg  confReg_6; // @[ScanConf.scala 32:20]
  reg  confReg_7; // @[ScanConf.scala 32:20]
  reg  confReg_8; // @[ScanConf.scala 32:20]
  reg  confReg_9; // @[ScanConf.scala 32:20]
  reg  confReg_10; // @[ScanConf.scala 32:20]
  reg  confReg_11; // @[ScanConf.scala 32:20]
  reg  confReg_12; // @[ScanConf.scala 32:20]
  reg  confReg_13; // @[ScanConf.scala 32:20]
  reg  confReg_14; // @[ScanConf.scala 32:20]
  reg  confReg_15; // @[ScanConf.scala 32:20]
  reg  confReg_16; // @[ScanConf.scala 32:20]
  reg  confReg_17; // @[ScanConf.scala 32:20]
  reg  confReg_18; // @[ScanConf.scala 32:20]
  reg  confReg_19; // @[ScanConf.scala 32:20]
  reg  confReg_20; // @[ScanConf.scala 32:20]
  reg  confReg_21; // @[ScanConf.scala 32:20]
  reg  confReg_22; // @[ScanConf.scala 32:20]
  reg  confReg_23; // @[ScanConf.scala 32:20]
  reg  confReg_24; // @[ScanConf.scala 32:20]
  reg  confReg_25; // @[ScanConf.scala 32:20]
  reg  confReg_26; // @[ScanConf.scala 32:20]
  reg  confReg_27; // @[ScanConf.scala 32:20]
  reg  confReg_28; // @[ScanConf.scala 32:20]
  reg  confReg_29; // @[ScanConf.scala 32:20]
  reg  confReg_30; // @[ScanConf.scala 32:20]
  reg  confReg_31; // @[ScanConf.scala 32:20]
  reg  confReg_32; // @[ScanConf.scala 32:20]
  reg  confReg_33; // @[ScanConf.scala 32:20]
  reg  confReg_34; // @[ScanConf.scala 32:20]
  reg  confReg_35; // @[ScanConf.scala 32:20]
  reg  confReg_36; // @[ScanConf.scala 32:20]
  reg  confReg_37; // @[ScanConf.scala 32:20]
  reg  confReg_38; // @[ScanConf.scala 32:20]
  reg  confReg_39; // @[ScanConf.scala 32:20]
  reg  confReg_40; // @[ScanConf.scala 32:20]
  reg  confReg_41; // @[ScanConf.scala 32:20]
  reg  confReg_42; // @[ScanConf.scala 32:20]
  reg  confReg_43; // @[ScanConf.scala 32:20]
  reg  confReg_44; // @[ScanConf.scala 32:20]
  reg  confReg_45; // @[ScanConf.scala 32:20]
  reg  confReg_46; // @[ScanConf.scala 32:20]
  reg  confReg_47; // @[ScanConf.scala 32:20]
  reg  confReg_48; // @[ScanConf.scala 32:20]
  reg  confReg_49; // @[ScanConf.scala 32:20]
  reg  confReg_50; // @[ScanConf.scala 32:20]
  reg  confReg_51; // @[ScanConf.scala 32:20]
  reg  confReg_52; // @[ScanConf.scala 32:20]
  reg  confReg_53; // @[ScanConf.scala 32:20]
  reg  confReg_54; // @[ScanConf.scala 32:20]
  reg  confReg_55; // @[ScanConf.scala 32:20]
  reg  confReg_56; // @[ScanConf.scala 32:20]
  reg  confReg_57; // @[ScanConf.scala 32:20]
  reg  confReg_58; // @[ScanConf.scala 32:20]
  reg  confReg_59; // @[ScanConf.scala 32:20]
  reg  confReg_60; // @[ScanConf.scala 32:20]
  reg  confReg_61; // @[ScanConf.scala 32:20]
  reg  confReg_62; // @[ScanConf.scala 32:20]
  reg  confReg_63; // @[ScanConf.scala 32:20]
  reg  confReg_64; // @[ScanConf.scala 32:20]
  reg  confReg_65; // @[ScanConf.scala 32:20]
  reg  confReg_66; // @[ScanConf.scala 32:20]
  reg  confReg_67; // @[ScanConf.scala 32:20]
  reg  confReg_68; // @[ScanConf.scala 32:20]
  reg  confReg_69; // @[ScanConf.scala 32:20]
  reg  confReg_70; // @[ScanConf.scala 32:20]
  reg  confReg_71; // @[ScanConf.scala 32:20]
  reg  confReg_72; // @[ScanConf.scala 32:20]
  reg  confReg_73; // @[ScanConf.scala 32:20]
  reg  confReg_74; // @[ScanConf.scala 32:20]
  reg  confReg_75; // @[ScanConf.scala 32:20]
  reg  confReg_76; // @[ScanConf.scala 32:20]
  reg  confReg_77; // @[ScanConf.scala 32:20]
  reg  confReg_78; // @[ScanConf.scala 32:20]
  reg  confReg_79; // @[ScanConf.scala 32:20]
  reg  confReg_80; // @[ScanConf.scala 32:20]
  reg  confReg_81; // @[ScanConf.scala 32:20]
  reg  confReg_82; // @[ScanConf.scala 32:20]
  reg  confReg_83; // @[ScanConf.scala 32:20]
  reg  confReg_84; // @[ScanConf.scala 32:20]
  reg  confReg_85; // @[ScanConf.scala 32:20]
  reg  confReg_86; // @[ScanConf.scala 32:20]
  reg  confReg_87; // @[ScanConf.scala 32:20]
  reg  confReg_88; // @[ScanConf.scala 32:20]
  reg  confReg_89; // @[ScanConf.scala 32:20]
  reg  confReg_90; // @[ScanConf.scala 32:20]
  reg  confReg_91; // @[ScanConf.scala 32:20]
  reg  confReg_92; // @[ScanConf.scala 32:20]
  reg  confReg_93; // @[ScanConf.scala 32:20]
  reg  confReg_94; // @[ScanConf.scala 32:20]
  reg  confReg_95; // @[ScanConf.scala 32:20]
  reg  confReg_96; // @[ScanConf.scala 32:20]
  reg  confReg_97; // @[ScanConf.scala 32:20]
  reg  confReg_98; // @[ScanConf.scala 32:20]
  reg  confReg_99; // @[ScanConf.scala 32:20]
  reg  confReg_100; // @[ScanConf.scala 32:20]
  reg  confReg_101; // @[ScanConf.scala 32:20]
  reg  confReg_102; // @[ScanConf.scala 32:20]
  reg  confReg_103; // @[ScanConf.scala 32:20]
  reg  confReg_104; // @[ScanConf.scala 32:20]
  reg  confReg_105; // @[ScanConf.scala 32:20]
  reg  confReg_106; // @[ScanConf.scala 32:20]
  reg  confReg_107; // @[ScanConf.scala 32:20]
  reg  confReg_108; // @[ScanConf.scala 32:20]
  reg  confReg_109; // @[ScanConf.scala 32:20]
  reg  confReg_110; // @[ScanConf.scala 32:20]
  reg  confReg_111; // @[ScanConf.scala 32:20]
  reg  confReg_112; // @[ScanConf.scala 32:20]
  reg  confReg_113; // @[ScanConf.scala 32:20]
  reg  confReg_114; // @[ScanConf.scala 32:20]
  reg  confReg_115; // @[ScanConf.scala 32:20]
  reg  confReg_116; // @[ScanConf.scala 32:20]
  reg  confReg_117; // @[ScanConf.scala 32:20]
  reg  confReg_118; // @[ScanConf.scala 32:20]
  reg  confReg_119; // @[ScanConf.scala 32:20]
  reg  confReg_120; // @[ScanConf.scala 32:20]
  reg  confReg_121; // @[ScanConf.scala 32:20]
  reg  confReg_122; // @[ScanConf.scala 32:20]
  reg  confReg_123; // @[ScanConf.scala 32:20]
  reg  confReg_124; // @[ScanConf.scala 32:20]
  reg  confReg_125; // @[ScanConf.scala 32:20]
  reg  confReg_126; // @[ScanConf.scala 32:20]
  reg  confReg_127; // @[ScanConf.scala 32:20]
  reg  confReg_128; // @[ScanConf.scala 32:20]
  reg  confReg_129; // @[ScanConf.scala 32:20]
  reg  confReg_130; // @[ScanConf.scala 32:20]
  reg  confReg_131; // @[ScanConf.scala 32:20]
  reg  confReg_132; // @[ScanConf.scala 32:20]
  reg  confReg_133; // @[ScanConf.scala 32:20]
  reg  confReg_134; // @[ScanConf.scala 32:20]
  reg  confReg_135; // @[ScanConf.scala 32:20]
  reg  confReg_136; // @[ScanConf.scala 32:20]
  reg  confReg_137; // @[ScanConf.scala 32:20]
  reg  confReg_138; // @[ScanConf.scala 32:20]
  reg  confReg_139; // @[ScanConf.scala 32:20]
  reg  confReg_140; // @[ScanConf.scala 32:20]
  reg  confReg_141; // @[ScanConf.scala 32:20]
  reg  confReg_142; // @[ScanConf.scala 32:20]
  reg  confReg_143; // @[ScanConf.scala 32:20]
  reg  confReg_144; // @[ScanConf.scala 32:20]
  reg  confReg_145; // @[ScanConf.scala 32:20]
  reg  confReg_146; // @[ScanConf.scala 32:20]
  reg  confReg_147; // @[ScanConf.scala 32:20]
  reg  confReg_148; // @[ScanConf.scala 32:20]
  reg  confReg_149; // @[ScanConf.scala 32:20]
  reg  confReg_150; // @[ScanConf.scala 32:20]
  reg  confReg_151; // @[ScanConf.scala 32:20]
  reg  confReg_152; // @[ScanConf.scala 32:20]
  reg  confReg_153; // @[ScanConf.scala 32:20]
  reg  confReg_154; // @[ScanConf.scala 32:20]
  reg  confReg_155; // @[ScanConf.scala 32:20]
  reg  confReg_156; // @[ScanConf.scala 32:20]
  reg  confReg_157; // @[ScanConf.scala 32:20]
  reg  confReg_158; // @[ScanConf.scala 32:20]
  reg  confReg_159; // @[ScanConf.scala 32:20]
  reg  confReg_160; // @[ScanConf.scala 32:20]
  reg  confReg_161; // @[ScanConf.scala 32:20]
  reg  confReg_162; // @[ScanConf.scala 32:20]
  reg  confReg_163; // @[ScanConf.scala 32:20]
  reg  confReg_164; // @[ScanConf.scala 32:20]
  reg  confReg_165; // @[ScanConf.scala 32:20]
  reg  confReg_166; // @[ScanConf.scala 32:20]
  reg  confReg_167; // @[ScanConf.scala 32:20]
  reg  confReg_168; // @[ScanConf.scala 32:20]
  reg  confReg_169; // @[ScanConf.scala 32:20]
  reg  confReg_170; // @[ScanConf.scala 32:20]
  reg  confReg_171; // @[ScanConf.scala 32:20]
  reg  confReg_172; // @[ScanConf.scala 32:20]
  reg  confReg_173; // @[ScanConf.scala 32:20]
  reg  confReg_174; // @[ScanConf.scala 32:20]
  reg  confReg_175; // @[ScanConf.scala 32:20]
  reg  confReg_176; // @[ScanConf.scala 32:20]
  reg  confReg_177; // @[ScanConf.scala 32:20]
  reg  confReg_178; // @[ScanConf.scala 32:20]
  reg  confReg_179; // @[ScanConf.scala 32:20]
  reg  confReg_180; // @[ScanConf.scala 32:20]
  reg  confReg_181; // @[ScanConf.scala 32:20]
  reg  confReg_182; // @[ScanConf.scala 32:20]
  reg  confReg_183; // @[ScanConf.scala 32:20]
  reg  confReg_184; // @[ScanConf.scala 32:20]
  reg  confReg_185; // @[ScanConf.scala 32:20]
  reg  confReg_186; // @[ScanConf.scala 32:20]
  reg  confReg_187; // @[ScanConf.scala 32:20]
  reg  confReg_188; // @[ScanConf.scala 32:20]
  reg  confReg_189; // @[ScanConf.scala 32:20]
  reg  confReg_190; // @[ScanConf.scala 32:20]
  reg  confReg_191; // @[ScanConf.scala 32:20]
  reg  confReg_192; // @[ScanConf.scala 32:20]
  reg  confReg_193; // @[ScanConf.scala 32:20]
  reg  confReg_194; // @[ScanConf.scala 32:20]
  reg  confReg_195; // @[ScanConf.scala 32:20]
  reg  confReg_196; // @[ScanConf.scala 32:20]
  reg  confReg_197; // @[ScanConf.scala 32:20]
  reg  confReg_198; // @[ScanConf.scala 32:20]
  reg  confReg_199; // @[ScanConf.scala 32:20]
  reg  confReg_200; // @[ScanConf.scala 32:20]
  reg  confReg_201; // @[ScanConf.scala 32:20]
  reg  confReg_202; // @[ScanConf.scala 32:20]
  reg  confReg_203; // @[ScanConf.scala 32:20]
  reg  confReg_204; // @[ScanConf.scala 32:20]
  reg  confReg_205; // @[ScanConf.scala 32:20]
  reg  confReg_206; // @[ScanConf.scala 32:20]
  reg  confReg_207; // @[ScanConf.scala 32:20]
  reg  confReg_208; // @[ScanConf.scala 32:20]
  reg  confReg_209; // @[ScanConf.scala 32:20]
  reg  confReg_210; // @[ScanConf.scala 32:20]
  reg  confReg_211; // @[ScanConf.scala 32:20]
  reg  confReg_212; // @[ScanConf.scala 32:20]
  reg  confReg_213; // @[ScanConf.scala 32:20]
  reg  confReg_214; // @[ScanConf.scala 32:20]
  reg  confReg_215; // @[ScanConf.scala 32:20]
  reg  confReg_216; // @[ScanConf.scala 32:20]
  reg  confReg_217; // @[ScanConf.scala 32:20]
  reg  confReg_218; // @[ScanConf.scala 32:20]
  reg  confReg_219; // @[ScanConf.scala 32:20]
  reg  confReg_220; // @[ScanConf.scala 32:20]
  reg  confReg_221; // @[ScanConf.scala 32:20]
  reg  confReg_222; // @[ScanConf.scala 32:20]
  reg  confReg_223; // @[ScanConf.scala 32:20]
  reg  confReg_224; // @[ScanConf.scala 32:20]
  reg  confReg_225; // @[ScanConf.scala 32:20]
  reg  confReg_226; // @[ScanConf.scala 32:20]
  reg  confReg_227; // @[ScanConf.scala 32:20]
  reg  confReg_228; // @[ScanConf.scala 32:20]
  reg  confReg_229; // @[ScanConf.scala 32:20]
  reg  confReg_230; // @[ScanConf.scala 32:20]
  reg  confReg_231; // @[ScanConf.scala 32:20]
  reg  confReg_232; // @[ScanConf.scala 32:20]
  reg  confReg_233; // @[ScanConf.scala 32:20]
  reg  confReg_234; // @[ScanConf.scala 32:20]
  reg  confReg_235; // @[ScanConf.scala 32:20]
  reg  confReg_236; // @[ScanConf.scala 32:20]
  reg  confReg_237; // @[ScanConf.scala 32:20]
  reg  confReg_238; // @[ScanConf.scala 32:20]
  reg  confReg_239; // @[ScanConf.scala 32:20]
  reg  confReg_240; // @[ScanConf.scala 32:20]
  reg  confReg_241; // @[ScanConf.scala 32:20]
  reg  confReg_242; // @[ScanConf.scala 32:20]
  reg  confReg_243; // @[ScanConf.scala 32:20]
  reg  confReg_244; // @[ScanConf.scala 32:20]
  reg  confReg_245; // @[ScanConf.scala 32:20]
  reg  confReg_246; // @[ScanConf.scala 32:20]
  reg  confReg_247; // @[ScanConf.scala 32:20]
  reg  confReg_248; // @[ScanConf.scala 32:20]
  reg  confReg_249; // @[ScanConf.scala 32:20]
  reg  confReg_250; // @[ScanConf.scala 32:20]
  reg  confReg_251; // @[ScanConf.scala 32:20]
  reg  confReg_252; // @[ScanConf.scala 32:20]
  reg  confReg_253; // @[ScanConf.scala 32:20]
  reg  confReg_254; // @[ScanConf.scala 32:20]
  reg  confReg_255; // @[ScanConf.scala 32:20]
  reg  confReg_256; // @[ScanConf.scala 32:20]
  reg  confReg_257; // @[ScanConf.scala 32:20]
  reg  confReg_258; // @[ScanConf.scala 32:20]
  reg  confReg_259; // @[ScanConf.scala 32:20]
  reg  confReg_260; // @[ScanConf.scala 32:20]
  reg  confReg_261; // @[ScanConf.scala 32:20]
  reg  confReg_262; // @[ScanConf.scala 32:20]
  reg  confReg_263; // @[ScanConf.scala 32:20]
  reg  confReg_264; // @[ScanConf.scala 32:20]
  reg  confReg_265; // @[ScanConf.scala 32:20]
  reg  confReg_266; // @[ScanConf.scala 32:20]
  reg  confReg_267; // @[ScanConf.scala 32:20]
  reg  confReg_268; // @[ScanConf.scala 32:20]
  reg  confReg_269; // @[ScanConf.scala 32:20]
  reg  confReg_270; // @[ScanConf.scala 32:20]
  reg  confReg_271; // @[ScanConf.scala 32:20]
  reg  confReg_272; // @[ScanConf.scala 32:20]
  reg  confReg_273; // @[ScanConf.scala 32:20]
  reg  confReg_274; // @[ScanConf.scala 32:20]
  reg  confReg_275; // @[ScanConf.scala 32:20]
  reg  confReg_276; // @[ScanConf.scala 32:20]
  reg  confReg_277; // @[ScanConf.scala 32:20]
  reg  confReg_278; // @[ScanConf.scala 32:20]
  reg  confReg_279; // @[ScanConf.scala 32:20]
  reg  confReg_280; // @[ScanConf.scala 32:20]
  reg  confReg_281; // @[ScanConf.scala 32:20]
  reg  confReg_282; // @[ScanConf.scala 32:20]
  reg  confReg_283; // @[ScanConf.scala 32:20]
  reg  confReg_284; // @[ScanConf.scala 32:20]
  reg  confReg_285; // @[ScanConf.scala 32:20]
  reg  confReg_286; // @[ScanConf.scala 32:20]
  reg  confReg_287; // @[ScanConf.scala 32:20]
  reg  confReg_288; // @[ScanConf.scala 32:20]
  reg  confReg_289; // @[ScanConf.scala 32:20]
  reg  confReg_290; // @[ScanConf.scala 32:20]
  reg  confReg_291; // @[ScanConf.scala 32:20]
  reg  confReg_292; // @[ScanConf.scala 32:20]
  reg  confReg_293; // @[ScanConf.scala 32:20]
  reg  confReg_294; // @[ScanConf.scala 32:20]
  reg  confReg_295; // @[ScanConf.scala 32:20]
  reg  confReg_296; // @[ScanConf.scala 32:20]
  reg  confReg_297; // @[ScanConf.scala 32:20]
  reg  confReg_298; // @[ScanConf.scala 32:20]
  reg  confReg_299; // @[ScanConf.scala 32:20]
  reg  confReg_300; // @[ScanConf.scala 32:20]
  reg  confReg_301; // @[ScanConf.scala 32:20]
  reg  confReg_302; // @[ScanConf.scala 32:20]
  reg  confReg_303; // @[ScanConf.scala 32:20]
  reg  confReg_304; // @[ScanConf.scala 32:20]
  reg  confReg_305; // @[ScanConf.scala 32:20]
  reg  confReg_306; // @[ScanConf.scala 32:20]
  reg  confReg_307; // @[ScanConf.scala 32:20]
  reg  confReg_308; // @[ScanConf.scala 32:20]
  reg  confReg_309; // @[ScanConf.scala 32:20]
  reg  confReg_310; // @[ScanConf.scala 32:20]
  reg  confReg_311; // @[ScanConf.scala 32:20]
  reg  confReg_312; // @[ScanConf.scala 32:20]
  reg  confReg_313; // @[ScanConf.scala 32:20]
  reg  confReg_314; // @[ScanConf.scala 32:20]
  reg  confReg_315; // @[ScanConf.scala 32:20]
  reg  confReg_316; // @[ScanConf.scala 32:20]
  reg  confReg_317; // @[ScanConf.scala 32:20]
  reg  confReg_318; // @[ScanConf.scala 32:20]
  reg  confReg_319; // @[ScanConf.scala 32:20]
  reg  confReg_320; // @[ScanConf.scala 32:20]
  reg  confReg_321; // @[ScanConf.scala 32:20]
  reg  confReg_322; // @[ScanConf.scala 32:20]
  reg  confReg_323; // @[ScanConf.scala 32:20]
  reg  confReg_324; // @[ScanConf.scala 32:20]
  reg  confReg_325; // @[ScanConf.scala 32:20]
  reg  confReg_326; // @[ScanConf.scala 32:20]
  reg  confReg_327; // @[ScanConf.scala 32:20]
  reg  confReg_328; // @[ScanConf.scala 32:20]
  reg  confReg_329; // @[ScanConf.scala 32:20]
  reg  confReg_330; // @[ScanConf.scala 32:20]
  reg  confReg_331; // @[ScanConf.scala 32:20]
  reg  confReg_332; // @[ScanConf.scala 32:20]
  reg  confReg_333; // @[ScanConf.scala 32:20]
  reg  confReg_334; // @[ScanConf.scala 32:20]
  reg  confReg_335; // @[ScanConf.scala 32:20]
  reg  confReg_336; // @[ScanConf.scala 32:20]
  reg  confReg_337; // @[ScanConf.scala 32:20]
  reg  confReg_338; // @[ScanConf.scala 32:20]
  reg  confReg_339; // @[ScanConf.scala 32:20]
  reg  confReg_340; // @[ScanConf.scala 32:20]
  reg  confReg_341; // @[ScanConf.scala 32:20]
  reg  confReg_342; // @[ScanConf.scala 32:20]
  reg  confReg_343; // @[ScanConf.scala 32:20]
  reg  confReg_344; // @[ScanConf.scala 32:20]
  reg  confReg_345; // @[ScanConf.scala 32:20]
  reg  confReg_346; // @[ScanConf.scala 32:20]
  reg  confReg_347; // @[ScanConf.scala 32:20]
  reg  confReg_348; // @[ScanConf.scala 32:20]
  reg  confReg_349; // @[ScanConf.scala 32:20]
  reg  confReg_350; // @[ScanConf.scala 32:20]
  reg  confReg_351; // @[ScanConf.scala 32:20]
  reg  confReg_352; // @[ScanConf.scala 32:20]
  reg  confReg_353; // @[ScanConf.scala 32:20]
  reg  confReg_354; // @[ScanConf.scala 32:20]
  reg  confReg_355; // @[ScanConf.scala 32:20]
  reg  confReg_356; // @[ScanConf.scala 32:20]
  reg  confReg_357; // @[ScanConf.scala 32:20]
  reg  confReg_358; // @[ScanConf.scala 32:20]
  reg  confReg_359; // @[ScanConf.scala 32:20]
  reg  confReg_360; // @[ScanConf.scala 32:20]
  reg  confReg_361; // @[ScanConf.scala 32:20]
  reg  confReg_362; // @[ScanConf.scala 32:20]
  reg  confReg_363; // @[ScanConf.scala 32:20]
  reg  confReg_364; // @[ScanConf.scala 32:20]
  reg  confReg_365; // @[ScanConf.scala 32:20]
  reg  confReg_366; // @[ScanConf.scala 32:20]
  reg  confReg_367; // @[ScanConf.scala 32:20]
  reg  confReg_368; // @[ScanConf.scala 32:20]
  reg  confReg_369; // @[ScanConf.scala 32:20]
  reg  confReg_370; // @[ScanConf.scala 32:20]
  reg  confReg_371; // @[ScanConf.scala 32:20]
  reg  confReg_372; // @[ScanConf.scala 32:20]
  reg  confReg_373; // @[ScanConf.scala 32:20]
  reg  confReg_374; // @[ScanConf.scala 32:20]
  reg  confReg_375; // @[ScanConf.scala 32:20]
  reg  confReg_376; // @[ScanConf.scala 32:20]
  reg  confReg_377; // @[ScanConf.scala 32:20]
  reg  confReg_378; // @[ScanConf.scala 32:20]
  reg  confReg_379; // @[ScanConf.scala 32:20]
  reg  confReg_380; // @[ScanConf.scala 32:20]
  reg  confReg_381; // @[ScanConf.scala 32:20]
  reg  confReg_382; // @[ScanConf.scala 32:20]
  reg  confReg_383; // @[ScanConf.scala 32:20]
  reg  confReg_384; // @[ScanConf.scala 32:20]
  reg  confReg_385; // @[ScanConf.scala 32:20]
  reg  confReg_386; // @[ScanConf.scala 32:20]
  reg  confReg_387; // @[ScanConf.scala 32:20]
  reg  confReg_388; // @[ScanConf.scala 32:20]
  reg  confReg_389; // @[ScanConf.scala 32:20]
  reg  confReg_390; // @[ScanConf.scala 32:20]
  reg  confReg_391; // @[ScanConf.scala 32:20]
  reg  confReg_392; // @[ScanConf.scala 32:20]
  reg  confReg_393; // @[ScanConf.scala 32:20]
  reg  confReg_394; // @[ScanConf.scala 32:20]
  reg  confReg_395; // @[ScanConf.scala 32:20]
  reg  confReg_396; // @[ScanConf.scala 32:20]
  reg  confReg_397; // @[ScanConf.scala 32:20]
  reg  confReg_398; // @[ScanConf.scala 32:20]
  reg  confReg_399; // @[ScanConf.scala 32:20]
  reg  confReg_400; // @[ScanConf.scala 32:20]
  reg  confReg_401; // @[ScanConf.scala 32:20]
  reg  confReg_402; // @[ScanConf.scala 32:20]
  reg  confReg_403; // @[ScanConf.scala 32:20]
  reg  confReg_404; // @[ScanConf.scala 32:20]
  reg  confReg_405; // @[ScanConf.scala 32:20]
  reg  confReg_406; // @[ScanConf.scala 32:20]
  reg  confReg_407; // @[ScanConf.scala 32:20]
  reg  confReg_408; // @[ScanConf.scala 32:20]
  reg  confReg_409; // @[ScanConf.scala 32:20]
  reg  confReg_410; // @[ScanConf.scala 32:20]
  reg  confReg_411; // @[ScanConf.scala 32:20]
  reg  confReg_412; // @[ScanConf.scala 32:20]
  reg  confReg_413; // @[ScanConf.scala 32:20]
  reg  confReg_414; // @[ScanConf.scala 32:20]
  reg  confReg_415; // @[ScanConf.scala 32:20]
  reg  confReg_416; // @[ScanConf.scala 32:20]
  reg  confReg_417; // @[ScanConf.scala 32:20]
  reg  confReg_418; // @[ScanConf.scala 32:20]
  reg  confReg_419; // @[ScanConf.scala 32:20]
  reg  confReg_420; // @[ScanConf.scala 32:20]
  reg  confReg_421; // @[ScanConf.scala 32:20]
  reg  confReg_422; // @[ScanConf.scala 32:20]
  reg  confReg_423; // @[ScanConf.scala 32:20]
  reg  confReg_424; // @[ScanConf.scala 32:20]
  reg  confReg_425; // @[ScanConf.scala 32:20]
  reg  confReg_426; // @[ScanConf.scala 32:20]
  reg  confReg_427; // @[ScanConf.scala 32:20]
  reg  confReg_428; // @[ScanConf.scala 32:20]
  reg  confReg_429; // @[ScanConf.scala 32:20]
  reg  confReg_430; // @[ScanConf.scala 32:20]
  reg  confReg_431; // @[ScanConf.scala 32:20]
  reg  confReg_432; // @[ScanConf.scala 32:20]
  reg  confReg_433; // @[ScanConf.scala 32:20]
  reg  confReg_434; // @[ScanConf.scala 32:20]
  reg  confReg_435; // @[ScanConf.scala 32:20]
  reg  confReg_436; // @[ScanConf.scala 32:20]
  reg  confReg_437; // @[ScanConf.scala 32:20]
  reg  confReg_438; // @[ScanConf.scala 32:20]
  reg  confReg_439; // @[ScanConf.scala 32:20]
  reg  confReg_440; // @[ScanConf.scala 32:20]
  reg  confReg_441; // @[ScanConf.scala 32:20]
  reg  confReg_442; // @[ScanConf.scala 32:20]
  reg  confReg_443; // @[ScanConf.scala 32:20]
  reg  confReg_444; // @[ScanConf.scala 32:20]
  reg  confReg_445; // @[ScanConf.scala 32:20]
  reg  confReg_446; // @[ScanConf.scala 32:20]
  reg  confReg_447; // @[ScanConf.scala 32:20]
  reg  confReg_448; // @[ScanConf.scala 32:20]
  reg  confReg_449; // @[ScanConf.scala 32:20]
  reg  confReg_450; // @[ScanConf.scala 32:20]
  reg  confReg_451; // @[ScanConf.scala 32:20]
  reg  confReg_452; // @[ScanConf.scala 32:20]
  reg  confReg_453; // @[ScanConf.scala 32:20]
  reg  confReg_454; // @[ScanConf.scala 32:20]
  reg  confReg_455; // @[ScanConf.scala 32:20]
  reg  confReg_456; // @[ScanConf.scala 32:20]
  reg  confReg_457; // @[ScanConf.scala 32:20]
  reg  confReg_458; // @[ScanConf.scala 32:20]
  reg  confReg_459; // @[ScanConf.scala 32:20]
  reg  confReg_460; // @[ScanConf.scala 32:20]
  reg  confReg_461; // @[ScanConf.scala 32:20]
  reg  confReg_462; // @[ScanConf.scala 32:20]
  reg  confReg_463; // @[ScanConf.scala 32:20]
  reg  confReg_464; // @[ScanConf.scala 32:20]
  reg  confReg_465; // @[ScanConf.scala 32:20]
  reg  confReg_466; // @[ScanConf.scala 32:20]
  reg  confReg_467; // @[ScanConf.scala 32:20]
  reg  confReg_468; // @[ScanConf.scala 32:20]
  reg  confReg_469; // @[ScanConf.scala 32:20]
  reg  confReg_470; // @[ScanConf.scala 32:20]
  reg  confReg_471; // @[ScanConf.scala 32:20]
  reg  confReg_472; // @[ScanConf.scala 32:20]
  reg  confReg_473; // @[ScanConf.scala 32:20]
  reg  confReg_474; // @[ScanConf.scala 32:20]
  reg  confReg_475; // @[ScanConf.scala 32:20]
  reg  confReg_476; // @[ScanConf.scala 32:20]
  reg  confReg_477; // @[ScanConf.scala 32:20]
  reg  confReg_478; // @[ScanConf.scala 32:20]
  reg  confReg_479; // @[ScanConf.scala 32:20]
  reg  confReg_480; // @[ScanConf.scala 32:20]
  reg  confReg_481; // @[ScanConf.scala 32:20]
  reg  confReg_482; // @[ScanConf.scala 32:20]
  reg  confReg_483; // @[ScanConf.scala 32:20]
  reg  confReg_484; // @[ScanConf.scala 32:20]
  reg  confReg_485; // @[ScanConf.scala 32:20]
  reg  confReg_486; // @[ScanConf.scala 32:20]
  reg  confReg_487; // @[ScanConf.scala 32:20]
  reg  confReg_488; // @[ScanConf.scala 32:20]
  reg  confReg_489; // @[ScanConf.scala 32:20]
  reg  confReg_490; // @[ScanConf.scala 32:20]
  reg  confReg_491; // @[ScanConf.scala 32:20]
  reg  confReg_492; // @[ScanConf.scala 32:20]
  reg  confReg_493; // @[ScanConf.scala 32:20]
  reg  confReg_494; // @[ScanConf.scala 32:20]
  reg  confReg_495; // @[ScanConf.scala 32:20]
  wire [3:0] io_scan_out_lo = {confReg_3,confReg_2,confReg_1,confReg_0}; // @[ScanConf.scala 46:47]
  wire [3:0] io_scan_out_hi = {confReg_7,confReg_6,confReg_5,confReg_4}; // @[ScanConf.scala 46:47]
  wire [6:0] io_confOut_lo_lo_lo_lo_lo_lo = {confReg_6,confReg_5,confReg_4,confReg_3,confReg_2,confReg_1,confReg_0}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_lo_lo_lo_lo_lo = {confReg_14,confReg_13,confReg_12,confReg_11,confReg_10,confReg_9,confReg_8,
    confReg_7,io_confOut_lo_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_lo_lo_hi_lo = {confReg_22,confReg_21,confReg_20,confReg_19,confReg_18,confReg_17,
    confReg_16,confReg_15}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_lo_lo_lo_lo = {confReg_30,confReg_29,confReg_28,confReg_27,confReg_26,confReg_25,confReg_24,
    confReg_23,io_confOut_lo_lo_lo_lo_hi_lo,io_confOut_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_lo_lo_hi_lo_lo = {confReg_37,confReg_36,confReg_35,confReg_34,confReg_33,confReg_32,
    confReg_31}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_lo_lo_lo_hi_lo = {confReg_45,confReg_44,confReg_43,confReg_42,confReg_41,confReg_40,confReg_39,
    confReg_38,io_confOut_lo_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_lo_hi_hi_lo = {confReg_53,confReg_52,confReg_51,confReg_50,confReg_49,confReg_48,
    confReg_47,confReg_46}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_lo_lo_lo_hi = {confReg_61,confReg_60,confReg_59,confReg_58,confReg_57,confReg_56,confReg_55,
    confReg_54,io_confOut_lo_lo_lo_hi_hi_lo,io_confOut_lo_lo_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_lo_hi_lo_lo_lo = {confReg_68,confReg_67,confReg_66,confReg_65,confReg_64,confReg_63,
    confReg_62}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_lo_lo_hi_lo_lo = {confReg_76,confReg_75,confReg_74,confReg_73,confReg_72,confReg_71,confReg_70,
    confReg_69,io_confOut_lo_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_hi_lo_hi_lo = {confReg_84,confReg_83,confReg_82,confReg_81,confReg_80,confReg_79,
    confReg_78,confReg_77}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_lo_lo_hi_lo = {confReg_92,confReg_91,confReg_90,confReg_89,confReg_88,confReg_87,confReg_86,
    confReg_85,io_confOut_lo_lo_hi_lo_hi_lo,io_confOut_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_lo_hi_hi_lo_lo = {confReg_99,confReg_98,confReg_97,confReg_96,confReg_95,confReg_94,
    confReg_93}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_lo_lo_hi_hi_lo = {confReg_107,confReg_106,confReg_105,confReg_104,confReg_103,confReg_102,
    confReg_101,confReg_100,io_confOut_lo_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_hi_hi_hi_lo = {confReg_115,confReg_114,confReg_113,confReg_112,confReg_111,confReg_110,
    confReg_109,confReg_108}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_lo_lo_hi_hi = {confReg_123,confReg_122,confReg_121,confReg_120,confReg_119,confReg_118,
    confReg_117,confReg_116,io_confOut_lo_lo_hi_hi_hi_lo,io_confOut_lo_lo_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_hi_lo_lo_lo_lo = {confReg_130,confReg_129,confReg_128,confReg_127,confReg_126,confReg_125,
    confReg_124}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_lo_hi_lo_lo_lo = {confReg_138,confReg_137,confReg_136,confReg_135,confReg_134,confReg_133,
    confReg_132,confReg_131,io_confOut_lo_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_lo_lo_hi_lo = {confReg_146,confReg_145,confReg_144,confReg_143,confReg_142,confReg_141,
    confReg_140,confReg_139}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_lo_hi_lo_lo = {confReg_154,confReg_153,confReg_152,confReg_151,confReg_150,confReg_149,
    confReg_148,confReg_147,io_confOut_lo_hi_lo_lo_hi_lo,io_confOut_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_hi_lo_hi_lo_lo = {confReg_161,confReg_160,confReg_159,confReg_158,confReg_157,confReg_156,
    confReg_155}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_lo_hi_lo_hi_lo = {confReg_169,confReg_168,confReg_167,confReg_166,confReg_165,confReg_164,
    confReg_163,confReg_162,io_confOut_lo_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_lo_hi_hi_lo = {confReg_177,confReg_176,confReg_175,confReg_174,confReg_173,confReg_172,
    confReg_171,confReg_170}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_lo_hi_lo_hi = {confReg_185,confReg_184,confReg_183,confReg_182,confReg_181,confReg_180,
    confReg_179,confReg_178,io_confOut_lo_hi_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_hi_hi_lo_lo_lo = {confReg_192,confReg_191,confReg_190,confReg_189,confReg_188,confReg_187,
    confReg_186}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_lo_hi_hi_lo_lo = {confReg_200,confReg_199,confReg_198,confReg_197,confReg_196,confReg_195,
    confReg_194,confReg_193,io_confOut_lo_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_hi_lo_hi_lo = {confReg_208,confReg_207,confReg_206,confReg_205,confReg_204,confReg_203,
    confReg_202,confReg_201}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_lo_hi_hi_lo = {confReg_216,confReg_215,confReg_214,confReg_213,confReg_212,confReg_211,
    confReg_210,confReg_209,io_confOut_lo_hi_hi_lo_hi_lo,io_confOut_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_lo_hi_hi_hi_lo_lo = {confReg_223,confReg_222,confReg_221,confReg_220,confReg_219,confReg_218,
    confReg_217}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_lo_hi_hi_hi_lo = {confReg_231,confReg_230,confReg_229,confReg_228,confReg_227,confReg_226,
    confReg_225,confReg_224,io_confOut_lo_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_hi_hi_hi_lo = {confReg_239,confReg_238,confReg_237,confReg_236,confReg_235,confReg_234,
    confReg_233,confReg_232}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_lo_hi_hi_hi = {confReg_247,confReg_246,confReg_245,confReg_244,confReg_243,confReg_242,
    confReg_241,confReg_240,io_confOut_lo_hi_hi_hi_hi_lo,io_confOut_lo_hi_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [247:0] io_confOut_lo = {io_confOut_lo_hi_hi_hi,io_confOut_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi,
    io_confOut_lo_hi_lo_lo,io_confOut_lo_lo_hi_hi,io_confOut_lo_lo_hi_lo,io_confOut_lo_lo_lo_hi,io_confOut_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_lo_lo_lo_lo_lo = {confReg_254,confReg_253,confReg_252,confReg_251,confReg_250,confReg_249,
    confReg_248}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_hi_lo_lo_lo_lo = {confReg_262,confReg_261,confReg_260,confReg_259,confReg_258,confReg_257,
    confReg_256,confReg_255,io_confOut_hi_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_lo_lo_hi_lo = {confReg_270,confReg_269,confReg_268,confReg_267,confReg_266,confReg_265,
    confReg_264,confReg_263}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_hi_lo_lo_lo = {confReg_278,confReg_277,confReg_276,confReg_275,confReg_274,confReg_273,
    confReg_272,confReg_271,io_confOut_hi_lo_lo_lo_hi_lo,io_confOut_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_lo_lo_hi_lo_lo = {confReg_285,confReg_284,confReg_283,confReg_282,confReg_281,confReg_280,
    confReg_279}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_hi_lo_lo_hi_lo = {confReg_293,confReg_292,confReg_291,confReg_290,confReg_289,confReg_288,
    confReg_287,confReg_286,io_confOut_hi_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_lo_hi_hi_lo = {confReg_301,confReg_300,confReg_299,confReg_298,confReg_297,confReg_296,
    confReg_295,confReg_294}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_hi_lo_lo_hi = {confReg_309,confReg_308,confReg_307,confReg_306,confReg_305,confReg_304,
    confReg_303,confReg_302,io_confOut_hi_lo_lo_hi_hi_lo,io_confOut_hi_lo_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_lo_hi_lo_lo_lo = {confReg_316,confReg_315,confReg_314,confReg_313,confReg_312,confReg_311,
    confReg_310}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_hi_lo_hi_lo_lo = {confReg_324,confReg_323,confReg_322,confReg_321,confReg_320,confReg_319,
    confReg_318,confReg_317,io_confOut_hi_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_hi_lo_hi_lo = {confReg_332,confReg_331,confReg_330,confReg_329,confReg_328,confReg_327,
    confReg_326,confReg_325}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_hi_lo_hi_lo = {confReg_340,confReg_339,confReg_338,confReg_337,confReg_336,confReg_335,
    confReg_334,confReg_333,io_confOut_hi_lo_hi_lo_hi_lo,io_confOut_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_lo_hi_hi_lo_lo = {confReg_347,confReg_346,confReg_345,confReg_344,confReg_343,confReg_342,
    confReg_341}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_hi_lo_hi_hi_lo = {confReg_355,confReg_354,confReg_353,confReg_352,confReg_351,confReg_350,
    confReg_349,confReg_348,io_confOut_hi_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_hi_hi_hi_lo = {confReg_363,confReg_362,confReg_361,confReg_360,confReg_359,confReg_358,
    confReg_357,confReg_356}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_hi_lo_hi_hi = {confReg_371,confReg_370,confReg_369,confReg_368,confReg_367,confReg_366,
    confReg_365,confReg_364,io_confOut_hi_lo_hi_hi_hi_lo,io_confOut_hi_lo_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_hi_lo_lo_lo_lo = {confReg_378,confReg_377,confReg_376,confReg_375,confReg_374,confReg_373,
    confReg_372}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_hi_hi_lo_lo_lo = {confReg_386,confReg_385,confReg_384,confReg_383,confReg_382,confReg_381,
    confReg_380,confReg_379,io_confOut_hi_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_lo_lo_hi_lo = {confReg_394,confReg_393,confReg_392,confReg_391,confReg_390,confReg_389,
    confReg_388,confReg_387}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_hi_hi_lo_lo = {confReg_402,confReg_401,confReg_400,confReg_399,confReg_398,confReg_397,
    confReg_396,confReg_395,io_confOut_hi_hi_lo_lo_hi_lo,io_confOut_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_hi_lo_hi_lo_lo = {confReg_409,confReg_408,confReg_407,confReg_406,confReg_405,confReg_404,
    confReg_403}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_hi_hi_lo_hi_lo = {confReg_417,confReg_416,confReg_415,confReg_414,confReg_413,confReg_412,
    confReg_411,confReg_410,io_confOut_hi_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_lo_hi_hi_lo = {confReg_425,confReg_424,confReg_423,confReg_422,confReg_421,confReg_420,
    confReg_419,confReg_418}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_hi_hi_lo_hi = {confReg_433,confReg_432,confReg_431,confReg_430,confReg_429,confReg_428,
    confReg_427,confReg_426,io_confOut_hi_hi_lo_hi_hi_lo,io_confOut_hi_hi_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_hi_hi_lo_lo_lo = {confReg_440,confReg_439,confReg_438,confReg_437,confReg_436,confReg_435,
    confReg_434}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_hi_hi_hi_lo_lo = {confReg_448,confReg_447,confReg_446,confReg_445,confReg_444,confReg_443,
    confReg_442,confReg_441,io_confOut_hi_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_hi_lo_hi_lo = {confReg_456,confReg_455,confReg_454,confReg_453,confReg_452,confReg_451,
    confReg_450,confReg_449}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_hi_hi_hi_lo = {confReg_464,confReg_463,confReg_462,confReg_461,confReg_460,confReg_459,
    confReg_458,confReg_457,io_confOut_hi_hi_hi_lo_hi_lo,io_confOut_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [6:0] io_confOut_hi_hi_hi_hi_lo_lo = {confReg_471,confReg_470,confReg_469,confReg_468,confReg_467,confReg_466,
    confReg_465}; // @[ScanConf.scala 48:25]
  wire [14:0] io_confOut_hi_hi_hi_hi_lo = {confReg_479,confReg_478,confReg_477,confReg_476,confReg_475,confReg_474,
    confReg_473,confReg_472,io_confOut_hi_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_hi_hi_hi_lo = {confReg_487,confReg_486,confReg_485,confReg_484,confReg_483,confReg_482,
    confReg_481,confReg_480}; // @[ScanConf.scala 48:25]
  wire [30:0] io_confOut_hi_hi_hi_hi = {confReg_495,confReg_494,confReg_493,confReg_492,confReg_491,confReg_490,
    confReg_489,confReg_488,io_confOut_hi_hi_hi_hi_hi_lo,io_confOut_hi_hi_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [247:0] io_confOut_hi = {io_confOut_hi_hi_hi_hi,io_confOut_hi_hi_hi_lo,io_confOut_hi_hi_lo_hi,
    io_confOut_hi_hi_lo_lo,io_confOut_hi_lo_hi_hi,io_confOut_hi_lo_hi_lo,io_confOut_hi_lo_lo_hi,io_confOut_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  assign ioBundle_confOut = {io_confOut_hi,io_confOut_lo}; // @[ScanConf.scala 48:25]
  assign ioBundle_scan_out = {io_scan_out_hi,io_scan_out_lo}; // @[ScanConf.scala 46:47]
  always @(posedge clock) begin
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_0 <= confReg_8; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_1 <= confReg_9; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_2 <= confReg_10; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_3 <= confReg_11; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_4 <= confReg_12; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_5 <= confReg_13; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_6 <= confReg_14; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_7 <= confReg_15; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_8 <= confReg_16; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_9 <= confReg_17; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_10 <= confReg_18; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_11 <= confReg_19; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_12 <= confReg_20; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_13 <= confReg_21; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_14 <= confReg_22; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_15 <= confReg_23; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_16 <= confReg_24; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_17 <= confReg_25; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_18 <= confReg_26; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_19 <= confReg_27; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_20 <= confReg_28; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_21 <= confReg_29; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_22 <= confReg_30; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_23 <= confReg_31; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_24 <= confReg_32; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_25 <= confReg_33; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_26 <= confReg_34; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_27 <= confReg_35; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_28 <= confReg_36; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_29 <= confReg_37; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_30 <= confReg_38; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_31 <= confReg_39; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_32 <= confReg_40; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_33 <= confReg_41; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_34 <= confReg_42; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_35 <= confReg_43; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_36 <= confReg_44; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_37 <= confReg_45; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_38 <= confReg_46; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_39 <= confReg_47; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_40 <= confReg_48; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_41 <= confReg_49; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_42 <= confReg_50; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_43 <= confReg_51; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_44 <= confReg_52; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_45 <= confReg_53; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_46 <= confReg_54; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_47 <= confReg_55; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_48 <= confReg_56; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_49 <= confReg_57; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_50 <= confReg_58; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_51 <= confReg_59; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_52 <= confReg_60; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_53 <= confReg_61; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_54 <= confReg_62; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_55 <= confReg_63; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_56 <= confReg_64; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_57 <= confReg_65; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_58 <= confReg_66; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_59 <= confReg_67; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_60 <= confReg_68; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_61 <= confReg_69; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_62 <= confReg_70; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_63 <= confReg_71; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_64 <= confReg_72; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_65 <= confReg_73; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_66 <= confReg_74; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_67 <= confReg_75; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_68 <= confReg_76; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_69 <= confReg_77; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_70 <= confReg_78; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_71 <= confReg_79; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_72 <= confReg_80; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_73 <= confReg_81; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_74 <= confReg_82; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_75 <= confReg_83; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_76 <= confReg_84; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_77 <= confReg_85; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_78 <= confReg_86; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_79 <= confReg_87; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_80 <= confReg_88; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_81 <= confReg_89; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_82 <= confReg_90; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_83 <= confReg_91; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_84 <= confReg_92; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_85 <= confReg_93; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_86 <= confReg_94; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_87 <= confReg_95; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_88 <= confReg_96; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_89 <= confReg_97; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_90 <= confReg_98; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_91 <= confReg_99; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_92 <= confReg_100; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_93 <= confReg_101; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_94 <= confReg_102; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_95 <= confReg_103; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_96 <= confReg_104; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_97 <= confReg_105; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_98 <= confReg_106; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_99 <= confReg_107; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_100 <= confReg_108; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_101 <= confReg_109; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_102 <= confReg_110; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_103 <= confReg_111; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_104 <= confReg_112; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_105 <= confReg_113; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_106 <= confReg_114; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_107 <= confReg_115; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_108 <= confReg_116; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_109 <= confReg_117; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_110 <= confReg_118; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_111 <= confReg_119; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_112 <= confReg_120; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_113 <= confReg_121; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_114 <= confReg_122; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_115 <= confReg_123; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_116 <= confReg_124; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_117 <= confReg_125; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_118 <= confReg_126; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_119 <= confReg_127; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_120 <= confReg_128; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_121 <= confReg_129; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_122 <= confReg_130; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_123 <= confReg_131; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_124 <= confReg_132; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_125 <= confReg_133; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_126 <= confReg_134; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_127 <= confReg_135; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_128 <= confReg_136; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_129 <= confReg_137; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_130 <= confReg_138; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_131 <= confReg_139; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_132 <= confReg_140; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_133 <= confReg_141; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_134 <= confReg_142; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_135 <= confReg_143; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_136 <= confReg_144; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_137 <= confReg_145; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_138 <= confReg_146; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_139 <= confReg_147; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_140 <= confReg_148; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_141 <= confReg_149; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_142 <= confReg_150; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_143 <= confReg_151; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_144 <= confReg_152; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_145 <= confReg_153; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_146 <= confReg_154; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_147 <= confReg_155; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_148 <= confReg_156; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_149 <= confReg_157; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_150 <= confReg_158; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_151 <= confReg_159; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_152 <= confReg_160; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_153 <= confReg_161; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_154 <= confReg_162; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_155 <= confReg_163; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_156 <= confReg_164; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_157 <= confReg_165; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_158 <= confReg_166; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_159 <= confReg_167; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_160 <= confReg_168; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_161 <= confReg_169; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_162 <= confReg_170; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_163 <= confReg_171; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_164 <= confReg_172; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_165 <= confReg_173; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_166 <= confReg_174; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_167 <= confReg_175; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_168 <= confReg_176; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_169 <= confReg_177; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_170 <= confReg_178; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_171 <= confReg_179; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_172 <= confReg_180; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_173 <= confReg_181; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_174 <= confReg_182; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_175 <= confReg_183; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_176 <= confReg_184; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_177 <= confReg_185; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_178 <= confReg_186; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_179 <= confReg_187; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_180 <= confReg_188; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_181 <= confReg_189; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_182 <= confReg_190; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_183 <= confReg_191; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_184 <= confReg_192; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_185 <= confReg_193; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_186 <= confReg_194; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_187 <= confReg_195; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_188 <= confReg_196; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_189 <= confReg_197; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_190 <= confReg_198; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_191 <= confReg_199; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_192 <= confReg_200; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_193 <= confReg_201; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_194 <= confReg_202; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_195 <= confReg_203; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_196 <= confReg_204; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_197 <= confReg_205; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_198 <= confReg_206; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_199 <= confReg_207; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_200 <= confReg_208; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_201 <= confReg_209; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_202 <= confReg_210; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_203 <= confReg_211; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_204 <= confReg_212; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_205 <= confReg_213; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_206 <= confReg_214; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_207 <= confReg_215; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_208 <= confReg_216; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_209 <= confReg_217; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_210 <= confReg_218; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_211 <= confReg_219; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_212 <= confReg_220; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_213 <= confReg_221; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_214 <= confReg_222; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_215 <= confReg_223; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_216 <= confReg_224; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_217 <= confReg_225; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_218 <= confReg_226; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_219 <= confReg_227; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_220 <= confReg_228; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_221 <= confReg_229; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_222 <= confReg_230; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_223 <= confReg_231; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_224 <= confReg_232; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_225 <= confReg_233; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_226 <= confReg_234; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_227 <= confReg_235; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_228 <= confReg_236; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_229 <= confReg_237; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_230 <= confReg_238; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_231 <= confReg_239; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_232 <= confReg_240; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_233 <= confReg_241; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_234 <= confReg_242; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_235 <= confReg_243; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_236 <= confReg_244; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_237 <= confReg_245; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_238 <= confReg_246; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_239 <= confReg_247; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_240 <= confReg_248; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_241 <= confReg_249; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_242 <= confReg_250; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_243 <= confReg_251; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_244 <= confReg_252; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_245 <= confReg_253; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_246 <= confReg_254; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_247 <= confReg_255; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_248 <= confReg_256; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_249 <= confReg_257; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_250 <= confReg_258; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_251 <= confReg_259; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_252 <= confReg_260; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_253 <= confReg_261; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_254 <= confReg_262; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_255 <= confReg_263; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_256 <= confReg_264; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_257 <= confReg_265; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_258 <= confReg_266; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_259 <= confReg_267; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_260 <= confReg_268; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_261 <= confReg_269; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_262 <= confReg_270; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_263 <= confReg_271; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_264 <= confReg_272; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_265 <= confReg_273; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_266 <= confReg_274; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_267 <= confReg_275; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_268 <= confReg_276; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_269 <= confReg_277; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_270 <= confReg_278; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_271 <= confReg_279; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_272 <= confReg_280; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_273 <= confReg_281; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_274 <= confReg_282; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_275 <= confReg_283; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_276 <= confReg_284; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_277 <= confReg_285; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_278 <= confReg_286; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_279 <= confReg_287; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_280 <= confReg_288; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_281 <= confReg_289; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_282 <= confReg_290; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_283 <= confReg_291; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_284 <= confReg_292; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_285 <= confReg_293; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_286 <= confReg_294; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_287 <= confReg_295; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_288 <= confReg_296; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_289 <= confReg_297; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_290 <= confReg_298; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_291 <= confReg_299; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_292 <= confReg_300; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_293 <= confReg_301; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_294 <= confReg_302; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_295 <= confReg_303; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_296 <= confReg_304; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_297 <= confReg_305; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_298 <= confReg_306; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_299 <= confReg_307; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_300 <= confReg_308; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_301 <= confReg_309; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_302 <= confReg_310; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_303 <= confReg_311; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_304 <= confReg_312; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_305 <= confReg_313; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_306 <= confReg_314; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_307 <= confReg_315; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_308 <= confReg_316; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_309 <= confReg_317; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_310 <= confReg_318; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_311 <= confReg_319; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_312 <= confReg_320; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_313 <= confReg_321; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_314 <= confReg_322; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_315 <= confReg_323; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_316 <= confReg_324; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_317 <= confReg_325; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_318 <= confReg_326; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_319 <= confReg_327; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_320 <= confReg_328; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_321 <= confReg_329; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_322 <= confReg_330; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_323 <= confReg_331; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_324 <= confReg_332; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_325 <= confReg_333; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_326 <= confReg_334; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_327 <= confReg_335; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_328 <= confReg_336; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_329 <= confReg_337; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_330 <= confReg_338; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_331 <= confReg_339; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_332 <= confReg_340; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_333 <= confReg_341; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_334 <= confReg_342; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_335 <= confReg_343; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_336 <= confReg_344; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_337 <= confReg_345; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_338 <= confReg_346; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_339 <= confReg_347; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_340 <= confReg_348; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_341 <= confReg_349; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_342 <= confReg_350; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_343 <= confReg_351; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_344 <= confReg_352; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_345 <= confReg_353; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_346 <= confReg_354; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_347 <= confReg_355; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_348 <= confReg_356; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_349 <= confReg_357; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_350 <= confReg_358; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_351 <= confReg_359; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_352 <= confReg_360; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_353 <= confReg_361; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_354 <= confReg_362; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_355 <= confReg_363; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_356 <= confReg_364; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_357 <= confReg_365; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_358 <= confReg_366; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_359 <= confReg_367; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_360 <= confReg_368; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_361 <= confReg_369; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_362 <= confReg_370; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_363 <= confReg_371; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_364 <= confReg_372; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_365 <= confReg_373; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_366 <= confReg_374; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_367 <= confReg_375; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_368 <= confReg_376; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_369 <= confReg_377; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_370 <= confReg_378; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_371 <= confReg_379; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_372 <= confReg_380; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_373 <= confReg_381; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_374 <= confReg_382; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_375 <= confReg_383; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_376 <= confReg_384; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_377 <= confReg_385; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_378 <= confReg_386; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_379 <= confReg_387; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_380 <= confReg_388; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_381 <= confReg_389; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_382 <= confReg_390; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_383 <= confReg_391; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_384 <= confReg_392; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_385 <= confReg_393; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_386 <= confReg_394; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_387 <= confReg_395; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_388 <= confReg_396; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_389 <= confReg_397; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_390 <= confReg_398; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_391 <= confReg_399; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_392 <= confReg_400; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_393 <= confReg_401; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_394 <= confReg_402; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_395 <= confReg_403; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_396 <= confReg_404; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_397 <= confReg_405; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_398 <= confReg_406; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_399 <= confReg_407; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_400 <= confReg_408; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_401 <= confReg_409; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_402 <= confReg_410; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_403 <= confReg_411; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_404 <= confReg_412; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_405 <= confReg_413; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_406 <= confReg_414; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_407 <= confReg_415; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_408 <= confReg_416; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_409 <= confReg_417; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_410 <= confReg_418; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_411 <= confReg_419; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_412 <= confReg_420; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_413 <= confReg_421; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_414 <= confReg_422; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_415 <= confReg_423; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_416 <= confReg_424; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_417 <= confReg_425; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_418 <= confReg_426; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_419 <= confReg_427; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_420 <= confReg_428; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_421 <= confReg_429; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_422 <= confReg_430; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_423 <= confReg_431; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_424 <= confReg_432; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_425 <= confReg_433; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_426 <= confReg_434; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_427 <= confReg_435; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_428 <= confReg_436; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_429 <= confReg_437; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_430 <= confReg_438; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_431 <= confReg_439; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_432 <= confReg_440; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_433 <= confReg_441; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_434 <= confReg_442; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_435 <= confReg_443; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_436 <= confReg_444; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_437 <= confReg_445; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_438 <= confReg_446; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_439 <= confReg_447; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_440 <= confReg_448; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_441 <= confReg_449; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_442 <= confReg_450; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_443 <= confReg_451; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_444 <= confReg_452; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_445 <= confReg_453; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_446 <= confReg_454; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_447 <= confReg_455; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_448 <= confReg_456; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_449 <= confReg_457; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_450 <= confReg_458; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_451 <= confReg_459; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_452 <= confReg_460; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_453 <= confReg_461; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_454 <= confReg_462; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_455 <= confReg_463; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_456 <= confReg_464; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_457 <= confReg_465; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_458 <= confReg_466; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_459 <= confReg_467; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_460 <= confReg_468; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_461 <= confReg_469; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_462 <= confReg_470; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_463 <= confReg_471; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_464 <= confReg_472; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_465 <= confReg_473; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_466 <= confReg_474; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_467 <= confReg_475; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_468 <= confReg_476; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_469 <= confReg_477; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_470 <= confReg_478; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_471 <= confReg_479; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_472 <= confReg_480; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_473 <= confReg_481; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_474 <= confReg_482; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_475 <= confReg_483; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_476 <= confReg_484; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_477 <= confReg_485; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_478 <= confReg_486; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_479 <= confReg_487; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_480 <= confReg_488; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_481 <= confReg_489; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_482 <= confReg_490; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_483 <= confReg_491; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_484 <= confReg_492; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_485 <= confReg_493; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_486 <= confReg_494; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_487 <= confReg_495; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_488 <= ioBundle_scan_in[0]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_489 <= ioBundle_scan_in[1]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_490 <= ioBundle_scan_in[2]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_491 <= ioBundle_scan_in[3]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_492 <= ioBundle_scan_in[4]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_493 <= ioBundle_scan_in[5]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_494 <= ioBundle_scan_in[6]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_495 <= ioBundle_scan_in[7]; // @[ScanConf.scala 38:72]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  confReg_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  confReg_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  confReg_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  confReg_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  confReg_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  confReg_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  confReg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  confReg_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  confReg_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  confReg_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  confReg_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  confReg_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  confReg_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  confReg_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  confReg_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  confReg_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  confReg_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  confReg_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  confReg_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  confReg_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  confReg_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  confReg_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  confReg_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  confReg_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  confReg_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  confReg_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  confReg_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  confReg_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  confReg_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  confReg_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  confReg_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  confReg_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  confReg_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  confReg_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  confReg_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  confReg_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  confReg_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  confReg_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  confReg_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  confReg_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  confReg_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  confReg_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  confReg_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  confReg_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  confReg_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  confReg_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  confReg_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  confReg_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  confReg_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  confReg_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  confReg_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  confReg_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  confReg_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  confReg_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  confReg_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  confReg_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  confReg_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  confReg_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  confReg_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  confReg_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  confReg_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  confReg_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  confReg_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  confReg_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  confReg_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  confReg_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  confReg_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  confReg_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  confReg_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  confReg_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  confReg_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  confReg_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  confReg_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  confReg_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  confReg_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  confReg_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  confReg_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  confReg_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  confReg_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  confReg_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  confReg_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  confReg_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  confReg_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  confReg_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  confReg_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  confReg_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  confReg_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  confReg_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  confReg_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  confReg_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  confReg_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  confReg_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  confReg_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  confReg_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  confReg_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  confReg_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  confReg_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  confReg_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  confReg_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  confReg_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  confReg_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  confReg_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  confReg_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  confReg_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  confReg_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  confReg_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  confReg_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  confReg_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  confReg_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  confReg_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  confReg_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  confReg_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  confReg_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  confReg_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  confReg_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  confReg_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  confReg_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  confReg_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  confReg_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  confReg_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  confReg_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  confReg_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  confReg_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  confReg_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  confReg_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  confReg_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  confReg_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  confReg_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  confReg_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  confReg_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  confReg_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  confReg_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  confReg_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  confReg_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  confReg_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  confReg_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  confReg_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  confReg_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  confReg_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  confReg_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  confReg_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  confReg_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  confReg_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  confReg_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  confReg_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  confReg_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  confReg_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  confReg_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  confReg_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  confReg_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  confReg_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  confReg_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  confReg_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  confReg_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  confReg_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  confReg_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  confReg_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  confReg_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  confReg_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  confReg_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  confReg_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  confReg_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  confReg_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  confReg_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  confReg_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  confReg_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  confReg_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  confReg_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  confReg_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  confReg_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  confReg_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  confReg_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  confReg_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  confReg_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  confReg_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  confReg_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  confReg_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  confReg_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  confReg_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  confReg_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  confReg_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  confReg_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  confReg_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  confReg_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  confReg_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  confReg_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  confReg_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  confReg_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  confReg_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  confReg_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  confReg_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  confReg_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  confReg_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  confReg_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  confReg_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  confReg_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  confReg_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  confReg_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  confReg_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  confReg_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  confReg_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  confReg_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  confReg_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  confReg_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  confReg_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  confReg_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  confReg_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  confReg_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  confReg_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  confReg_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  confReg_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  confReg_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  confReg_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  confReg_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  confReg_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  confReg_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  confReg_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  confReg_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  confReg_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  confReg_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  confReg_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  confReg_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  confReg_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  confReg_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  confReg_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  confReg_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  confReg_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  confReg_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  confReg_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  confReg_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  confReg_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  confReg_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  confReg_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  confReg_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  confReg_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  confReg_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  confReg_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  confReg_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  confReg_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  confReg_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  confReg_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  confReg_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  confReg_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  confReg_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  confReg_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  confReg_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  confReg_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  confReg_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  confReg_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  confReg_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  confReg_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  confReg_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  confReg_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  confReg_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  confReg_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  confReg_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  confReg_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  confReg_257 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  confReg_258 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  confReg_259 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  confReg_260 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  confReg_261 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  confReg_262 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  confReg_263 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  confReg_264 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  confReg_265 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  confReg_266 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  confReg_267 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  confReg_268 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  confReg_269 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  confReg_270 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  confReg_271 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  confReg_272 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  confReg_273 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  confReg_274 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  confReg_275 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  confReg_276 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  confReg_277 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  confReg_278 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  confReg_279 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  confReg_280 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  confReg_281 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  confReg_282 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  confReg_283 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  confReg_284 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  confReg_285 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  confReg_286 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  confReg_287 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  confReg_288 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  confReg_289 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  confReg_290 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  confReg_291 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  confReg_292 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  confReg_293 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  confReg_294 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  confReg_295 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  confReg_296 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  confReg_297 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  confReg_298 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  confReg_299 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  confReg_300 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  confReg_301 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  confReg_302 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  confReg_303 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  confReg_304 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  confReg_305 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  confReg_306 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  confReg_307 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  confReg_308 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  confReg_309 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  confReg_310 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  confReg_311 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  confReg_312 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  confReg_313 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  confReg_314 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  confReg_315 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  confReg_316 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  confReg_317 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  confReg_318 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  confReg_319 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  confReg_320 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  confReg_321 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  confReg_322 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  confReg_323 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  confReg_324 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  confReg_325 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  confReg_326 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  confReg_327 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  confReg_328 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  confReg_329 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  confReg_330 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  confReg_331 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  confReg_332 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  confReg_333 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  confReg_334 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  confReg_335 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  confReg_336 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  confReg_337 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  confReg_338 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  confReg_339 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  confReg_340 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  confReg_341 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  confReg_342 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  confReg_343 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  confReg_344 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  confReg_345 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  confReg_346 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  confReg_347 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  confReg_348 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  confReg_349 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  confReg_350 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  confReg_351 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  confReg_352 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  confReg_353 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  confReg_354 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  confReg_355 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  confReg_356 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  confReg_357 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  confReg_358 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  confReg_359 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  confReg_360 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  confReg_361 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  confReg_362 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  confReg_363 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  confReg_364 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  confReg_365 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  confReg_366 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  confReg_367 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  confReg_368 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  confReg_369 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  confReg_370 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  confReg_371 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  confReg_372 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  confReg_373 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  confReg_374 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  confReg_375 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  confReg_376 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  confReg_377 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  confReg_378 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  confReg_379 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  confReg_380 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  confReg_381 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  confReg_382 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  confReg_383 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  confReg_384 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  confReg_385 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  confReg_386 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  confReg_387 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  confReg_388 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  confReg_389 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  confReg_390 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  confReg_391 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  confReg_392 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  confReg_393 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  confReg_394 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  confReg_395 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  confReg_396 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  confReg_397 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  confReg_398 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  confReg_399 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  confReg_400 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  confReg_401 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  confReg_402 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  confReg_403 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  confReg_404 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  confReg_405 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  confReg_406 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  confReg_407 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  confReg_408 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  confReg_409 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  confReg_410 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  confReg_411 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  confReg_412 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  confReg_413 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  confReg_414 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  confReg_415 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  confReg_416 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  confReg_417 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  confReg_418 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  confReg_419 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  confReg_420 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  confReg_421 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  confReg_422 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  confReg_423 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  confReg_424 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  confReg_425 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  confReg_426 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  confReg_427 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  confReg_428 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  confReg_429 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  confReg_430 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  confReg_431 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  confReg_432 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  confReg_433 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  confReg_434 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  confReg_435 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  confReg_436 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  confReg_437 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  confReg_438 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  confReg_439 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  confReg_440 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  confReg_441 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  confReg_442 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  confReg_443 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  confReg_444 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  confReg_445 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  confReg_446 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  confReg_447 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  confReg_448 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  confReg_449 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  confReg_450 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  confReg_451 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  confReg_452 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  confReg_453 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  confReg_454 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  confReg_455 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  confReg_456 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  confReg_457 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  confReg_458 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  confReg_459 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  confReg_460 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  confReg_461 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  confReg_462 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  confReg_463 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  confReg_464 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  confReg_465 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  confReg_466 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  confReg_467 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  confReg_468 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  confReg_469 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  confReg_470 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  confReg_471 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  confReg_472 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  confReg_473 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  confReg_474 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  confReg_475 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  confReg_476 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  confReg_477 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  confReg_478 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  confReg_479 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  confReg_480 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  confReg_481 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  confReg_482 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  confReg_483 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  confReg_484 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  confReg_485 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  confReg_486 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  confReg_487 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  confReg_488 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  confReg_489 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  confReg_490 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  confReg_491 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  confReg_492 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  confReg_493 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  confReg_494 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  confReg_495 = _RAND_495[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MuxNInput_10_SCAOptCB(
  input  [9:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_cnstClk,
  input        io_arst
);
  wire [15:0] OPinMux_in; // @[MuxListTest.scala 43:28]
  wire [3:0] OPinMux_sel; // @[MuxListTest.scala 43:28]
  wire  OPinMux_o; // @[MuxListTest.scala 43:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux16C OPinMux ( // @[MuxListTest.scala 43:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{6'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_12_SCAOptCB(
  input  [11:0] io_in,
  input  [3:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [15:0] OPinMux_in; // @[MuxListTest.scala 43:28]
  wire [3:0] OPinMux_sel; // @[MuxListTest.scala 43:28]
  wire  OPinMux_o; // @[MuxListTest.scala 43:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux16C OPinMux ( // @[MuxListTest.scala 43:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{4'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_14_SCAOptCB(
  input  [13:0] io_in,
  input  [3:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [15:0] OPinMux_in; // @[MuxListTest.scala 43:28]
  wire [3:0] OPinMux_sel; // @[MuxListTest.scala 43:28]
  wire  OPinMux_o; // @[MuxListTest.scala 43:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux16C OPinMux ( // @[MuxListTest.scala 43:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{2'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_8_SCAOptCB(
  input  [7:0] io_in,
  input  [3:0] io_config,
  input        io_loopBreak,
  input        io_cnstClk,
  input        io_arst
);
  wire [15:0] OPinMux_in; // @[MuxListTest.scala 43:28]
  wire [3:0] OPinMux_sel; // @[MuxListTest.scala 43:28]
  wire  OPinMux_o; // @[MuxListTest.scala 43:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux16C OPinMux ( // @[MuxListTest.scala 43:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign OPinMux_in = {{8'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_O3_C6_SCAOptSB(
  input  [8:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{5'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in[8:3]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O3_C5_SCAOptSB(
  input  [7:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{5'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in[7:3]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O0_C6_SCAOptSB(
  input  [5:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = 8'h0; // @[MuxListTest.scala 125:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O0_C4_SCAOptSB(
  input  [3:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = 4'h0; // @[MuxListTest.scala 125:22]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = io_in; // @[MuxListTest.scala 144:28]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O4_C6_SCAOptSB(
  input  [9:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{4'd0}, io_in[3:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in[9:4]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O4_C5_SCAOptSB(
  input  [8:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{4'd0}, io_in[3:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in[8:4]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O4_C7_SCAOptSB(
  input  [10:0] io_in,
  input  [3:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_ioGndBle,
  input         io_cnstClk,
  input         io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{4'd0}, io_in[3:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{1'd0}, io_in[10:4]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module MuxNInput_O3_C7_SCAOptSB(
  input  [9:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 148:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 148:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 149:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 149:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 148:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 149:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 157:25]
  assign OPinMux_in = {{5'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{1'd0}, io_in[9:3]}; // @[MuxListTest.scala 144:20]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 155:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 156:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 154:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 150:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 152:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 151:17]
endmodule
module Tile_9_3_clbmemtile(
  input          clock,
  input          reset,
  input          IN_OPIN_N19967_41,
  input          IN_OPIN_N19968_42,
  input          IN_OPIN_N19969_43,
  input          IN_OPIN_N19970_44,
  input          IN_OPIN_N19971_45,
  input          IN_OPIN_N19972_46,
  input          IN_OPIN_N19973_47,
  input          IN_OPIN_N19974_48,
  input          IN_OPIN_N21019_49,
  input          IN_OPIN_N21020_50,
  input          IN_OPIN_N21021_51,
  input          IN_OPIN_N21022_52,
  input          IN_OPIN_N21023_53,
  input          IN_OPIN_N21024_54,
  input          IN_OPIN_N21025_55,
  input          IN_OPIN_N21026_56,
  input          IN_CHANX_N24152_0,
  input          IN_CHANX_N24154_8,
  input          IN_CHANX_N24156_16,
  input          IN_CHANX_N24158_24,
  input          IN_CHANX_N24160_32,
  input          IN_CHANX_N24162_40,
  input          IN_CHANX_N24164_48,
  input          IN_CHANX_N24166_56,
  input          IN_CHANX_N24168_64,
  input          IN_CHANX_N24170_72,
  input          IN_CHANX_N24174_2,
  input          IN_CHANX_N24175_3,
  input          IN_CHANX_N24176_10,
  input          IN_CHANX_N24177_11,
  input          IN_CHANX_N24178_18,
  input          IN_CHANX_N24179_19,
  input          IN_CHANX_N24180_26,
  input          IN_CHANX_N24181_27,
  input          IN_CHANX_N24182_34,
  input          IN_CHANX_N24183_35,
  input          IN_CHANX_N24196_4,
  input          IN_CHANX_N24197_5,
  input          IN_CHANX_N24198_12,
  input          IN_CHANX_N24199_13,
  input          IN_CHANX_N24200_20,
  input          IN_CHANX_N24201_21,
  input          IN_CHANX_N24202_28,
  input          IN_CHANX_N24203_29,
  input          IN_CHANX_N24204_36,
  input          IN_CHANX_N24205_37,
  input          IN_CHANX_N24214_76,
  input          IN_CHANX_N24216_6,
  input          IN_CHANX_N24217_7,
  input          IN_CHANX_N24218_14,
  input          IN_CHANX_N24219_15,
  input          IN_CHANX_N24220_22,
  input          IN_CHANX_N24221_23,
  input          IN_CHANX_N24222_30,
  input          IN_CHANX_N24223_31,
  input          IN_CHANX_N24224_38,
  input          IN_CHANX_N24225_39,
  input          IN_CHANX_N24226_46,
  input          IN_CHANX_N24227_47,
  input          IN_CHANX_N24228_54,
  input          IN_CHANX_N24229_55,
  input          IN_CHANX_N24230_62,
  input          IN_CHANX_N24231_63,
  input          IN_CHANX_N24232_70,
  input          IN_CHANX_N24233_71,
  input          IN_CHANX_N24237_1,
  input          IN_CHANX_N24239_9,
  input          IN_CHANX_N24241_17,
  input          IN_CHANX_N24243_25,
  input          IN_CHANX_N24245_33,
  input          IN_CHANX_N24247_41,
  input          IN_CHANX_N24249_49,
  input          IN_CHANX_N24251_57,
  input          IN_CHANX_N24253_65,
  input          IN_CHANX_N24255_73,
  input          IN_CHANX_N24257_77,
  input          IN_CHANY_N28730_0,
  input          IN_CHANY_N28732_2,
  input          IN_CHANY_N28733_3,
  input          IN_CHANY_N28738_8,
  input          IN_CHANY_N28740_10,
  input          IN_CHANY_N28741_11,
  input          IN_CHANY_N28746_16,
  input          IN_CHANY_N28748_18,
  input          IN_CHANY_N28749_19,
  input          IN_CHANY_N28754_24,
  input          IN_CHANY_N28756_26,
  input          IN_CHANY_N28757_27,
  input          IN_CHANY_N28762_32,
  input          IN_CHANY_N28764_34,
  input          IN_CHANY_N28765_35,
  input          IN_CHANY_N28770_40,
  input          IN_CHANY_N28778_48,
  input          IN_CHANY_N28786_56,
  input          IN_CHANY_N28794_64,
  input          IN_CHANY_N28802_72,
  input          IN_CHANY_N28810_4,
  input          IN_CHANY_N28811_5,
  input          IN_CHANY_N28812_12,
  input          IN_CHANY_N28813_13,
  input          IN_CHANY_N28814_20,
  input          IN_CHANY_N28815_21,
  input          IN_CHANY_N28816_28,
  input          IN_CHANY_N28817_29,
  input          IN_CHANY_N28818_36,
  input          IN_CHANY_N28819_37,
  input          IN_CHANY_N28828_76,
  input          IN_CHANY_N28830_6,
  input          IN_CHANY_N28831_7,
  input          IN_CHANY_N28832_14,
  input          IN_CHANY_N28833_15,
  input          IN_CHANY_N28834_22,
  input          IN_CHANY_N28835_23,
  input          IN_CHANY_N28836_30,
  input          IN_CHANY_N28837_31,
  input          IN_CHANY_N28838_38,
  input          IN_CHANY_N28839_39,
  input          IN_CHANY_N28840_46,
  input          IN_CHANY_N28841_47,
  input          IN_CHANY_N28842_54,
  input          IN_CHANY_N28843_55,
  input          IN_CHANY_N28844_62,
  input          IN_CHANY_N28845_63,
  input          IN_CHANY_N28846_70,
  input          IN_CHANY_N28847_71,
  input          IN_CHANY_N28848_78,
  input          IN_CHANY_N28849_79,
  input          IN_CHANY_N28851_1,
  input          IN_CHANY_N28853_9,
  input          IN_CHANY_N28855_17,
  input          IN_CHANY_N28857_25,
  input          IN_CHANY_N28859_33,
  input          IN_CHANY_N28861_41,
  input          IN_CHANY_N28863_49,
  input          IN_CHANY_N28865_57,
  input          IN_CHANY_N28867_65,
  input          IN_CHANY_N28869_73,
  input          IN_CHANY_N28871_77,
  output         OUT_CHANX_N24242_24,
  output         OUT_CHANX_N24250_56,
  output         OUT_CHANX_N24159_25,
  output         OUT_CHANY_N28868_72,
  output         OUT_CHANY_N28771_41,
  output         OUT_CHANY_N28747_17,
  output         OUT_CHANY_N28858_32,
  output         OUT_OPIN_N19855_45,
  output         OUT_CHANY_N28866_64,
  output         OUT_CHANY_N28829_77,
  output         OUT_OPIN_N19861_51,
  output         OUT_CHANX_N24171_73,
  output         OUT_CHANX_N24155_9,
  output         OUT_CHANX_N24161_33,
  output         OUT_CHANX_N24246_40,
  output         OUT_CHANX_N24165_49,
  output         OUT_CHANX_N24153_1,
  output         OUT_OPIN_N19860_50,
  output         OUT_CHANX_N24244_32,
  output         OUT_OPIN_N19858_48,
  output         OUT_CHANX_N24163_41,
  output         OUT_CHANY_N28739_9,
  output         OUT_OPIN_N19864_54,
  output         OUT_CHANY_N28860_40,
  output         OUT_CHANY_N28864_56,
  output         OUT_CHANY_N28850_0,
  output         OUT_CHANY_N28755_25,
  output         OUT_CHANY_N28731_1,
  output         OUT_OPIN_N19865_55,
  output         OUT_CHANX_N24252_64,
  output         OUT_CHANY_N28870_76,
  output         OUT_CHANY_N28795_65,
  output         OUT_CHANY_N28856_24,
  output         OUT_CHANX_N24240_16,
  output         OUT_CHANX_N24238_8,
  output         OUT_OPIN_N19854_44,
  output         OUT_CHANY_N28862_48,
  output         OUT_OPIN_N19851_41,
  output         OUT_CHANX_N24215_77,
  output         OUT_CHANX_N24256_76,
  output         OUT_OPIN_N19853_43,
  output         OUT_CHANX_N24254_72,
  output         OUT_CHANX_N24248_48,
  output         OUT_OPIN_N19857_47,
  output         OUT_CHANY_N28779_49,
  output         OUT_OPIN_N19856_46,
  output         OUT_CHANX_N24236_0,
  output         OUT_OPIN_N19863_53,
  output         OUT_CHANY_N28854_16,
  output         OUT_OPIN_N19859_49,
  output         OUT_CHANY_N28803_73,
  output         OUT_CHANX_N24167_57,
  output         OUT_OPIN_N19866_56,
  output         OUT_OPIN_N19852_42,
  output         OUT_CHANY_N28763_33,
  output         OUT_CHANX_N24157_17,
  output         OUT_CHANY_N28852_8,
  output         OUT_CHANX_N24169_65,
  output         OUT_CHANY_N28787_57,
  output         OUT_OPIN_N19862_52,
  output [495:0] ioConf_confOut,
  input  [7:0]   ioConf_scan_in,
  input          ioConf_scan_en,
  output [7:0]   ioConf_scan_out,
  input  [31:0]  ioPad_i,
  input          ctrlSignals_gndBlkOuts,
  input          ctrlSignals_loopBreak,
  input          ctrlSignals_arst,
  input          ctrlSignals_tmrMode,
  input          ctrlSignals_confClock,
  input          ctrlSignals_constClock
);
  wire  logicBlock_IPIN_0; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_1; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_2; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_3; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_4; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_5; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_6; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_7; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_8; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_9; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_10; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_11; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_12; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_13; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_14; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_15; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_16; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_17; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_18; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_19; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_20; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_21; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_22; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_23; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_24; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_25; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_26; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_27; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_28; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_29; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_30; // @[TileFull.scala 46:37]
  wire  logicBlock_IPIN_31; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_41; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_42; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_43; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_44; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_45; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_46; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_47; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_48; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_49; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_50; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_51; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_52; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_53; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_54; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_55; // @[TileFull.scala 46:37]
  wire  logicBlock_OPIN_56; // @[TileFull.scala 46:37]
  wire  logicBlock_clock; // @[TileFull.scala 46:37]
  wire  logicBlock_reset; // @[TileFull.scala 46:37]
  wire [15:0] logicBlock_ioPad_i; // @[TileFull.scala 46:37]
  wire [161:0] logicBlock_configBits; // @[TileFull.scala 46:37]
  wire  logicBlock_gndLBouts; // @[TileFull.scala 46:37]
  wire  configBlock_clock; // @[TileFull.scala 61:31]
  wire [495:0] configBlock_ioBundle_confOut; // @[TileFull.scala 61:31]
  wire [7:0] configBlock_ioBundle_scan_in; // @[TileFull.scala 61:31]
  wire  configBlock_ioBundle_scan_en; // @[TileFull.scala 61:31]
  wire [7:0] configBlock_ioBundle_scan_out; // @[TileFull.scala 61:31]
  wire [9:0] CBMux_IPIN0_N19810_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN0_N19810_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N19810_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N19810_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N19810_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN0_N19810_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN1_N19811_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN1_N19811_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN1_N19811_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN1_N19811_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN1_N19811_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN1_N19811_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN2_N19812_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN2_N19812_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N19812_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N19812_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N19812_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN2_N19812_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN3_N19813_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN3_N19813_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN3_N19813_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN3_N19813_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN3_N19813_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN3_N19813_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN4_N19814_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN4_N19814_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N19814_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N19814_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N19814_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN4_N19814_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN5_N19815_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN5_N19815_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN5_N19815_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN5_N19815_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN5_N19815_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN5_N19815_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN6_N19816_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN6_N19816_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N19816_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N19816_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N19816_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN6_N19816_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN7_N19817_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN7_N19817_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN7_N19817_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN7_N19817_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN7_N19817_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN7_N19817_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN8_N19818_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN8_N19818_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N19818_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N19818_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N19818_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN8_N19818_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN9_N19819_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN9_N19819_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN9_N19819_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN9_N19819_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN9_N19819_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN9_N19819_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN10_N19820_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN10_N19820_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N19820_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N19820_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N19820_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN10_N19820_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN11_N19821_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN11_N19821_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN11_N19821_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN11_N19821_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN11_N19821_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN11_N19821_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN12_N19822_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN12_N19822_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N19822_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N19822_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N19822_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN12_N19822_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN13_N19823_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN13_N19823_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN13_N19823_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN13_N19823_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN13_N19823_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN13_N19823_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN14_N19824_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN14_N19824_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N19824_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N19824_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N19824_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN14_N19824_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN15_N19825_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN15_N19825_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN15_N19825_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN15_N19825_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN15_N19825_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN15_N19825_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN16_N19826_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN16_N19826_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N19826_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N19826_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N19826_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN16_N19826_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN17_N19827_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN17_N19827_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN17_N19827_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN17_N19827_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN17_N19827_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN17_N19827_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN18_N19828_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN18_N19828_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N19828_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N19828_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N19828_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN18_N19828_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN19_N19829_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN19_N19829_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN19_N19829_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN19_N19829_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN19_N19829_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN19_N19829_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN20_N19830_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN20_N19830_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N19830_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N19830_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N19830_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN20_N19830_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN21_N19831_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN21_N19831_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN21_N19831_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN21_N19831_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN21_N19831_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN21_N19831_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN22_N19832_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN22_N19832_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N19832_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N19832_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N19832_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN22_N19832_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN23_N19833_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN23_N19833_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN23_N19833_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN23_N19833_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN23_N19833_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN23_N19833_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN24_N19834_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN24_N19834_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N19834_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N19834_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N19834_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN24_N19834_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN25_N19835_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN25_N19835_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN25_N19835_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN25_N19835_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN25_N19835_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN25_N19835_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN26_N19836_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN26_N19836_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N19836_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N19836_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N19836_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN26_N19836_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN27_N19837_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN27_N19837_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN27_N19837_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN27_N19837_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN27_N19837_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN27_N19837_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN28_N19838_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN28_N19838_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N19838_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N19838_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N19838_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN28_N19838_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN29_N19839_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN29_N19839_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN29_N19839_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN29_N19839_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN29_N19839_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN29_N19839_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN30_N19840_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN30_N19840_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N19840_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N19840_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N19840_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN30_N19840_io_arst; // @[TileFull.scala 97:27]
  wire [13:0] CBMux_IPIN31_N19841_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN31_N19841_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN31_N19841_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN31_N19841_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN31_N19841_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN31_N19841_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN32_N19842_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN32_N19842_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N19842_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N19842_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N19842_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN32_N19842_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN33_N19843_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN33_N19843_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN33_N19843_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN33_N19843_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN33_N19843_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN33_N19843_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN34_N19844_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN34_N19844_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N19844_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N19844_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N19844_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN34_N19844_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN35_N19845_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN35_N19845_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN35_N19845_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN35_N19845_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN35_N19845_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN35_N19845_io_arst; // @[TileFull.scala 97:27]
  wire [7:0] CBMux_IPIN36_N19846_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN36_N19846_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N19846_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N19846_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN36_N19846_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN37_N19847_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN37_N19847_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN37_N19847_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN37_N19847_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN37_N19847_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN37_N19847_io_arst; // @[TileFull.scala 97:27]
  wire [11:0] CBMux_IPIN38_N19848_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN38_N19848_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N19848_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N19848_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N19848_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN38_N19848_io_arst; // @[TileFull.scala 97:27]
  wire [9:0] CBMux_IPIN39_N19849_io_in; // @[TileFull.scala 97:27]
  wire [3:0] CBMux_IPIN39_N19849_io_config; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN39_N19849_io_out; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN39_N19849_io_loopBreak; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN39_N19849_io_cnstClk; // @[TileFull.scala 97:27]
  wire  CBMux_IPIN39_N19849_io_arst; // @[TileFull.scala 97:27]
  wire [8:0] SBMux_C1_N24153_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C1_N24153_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N24153_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N24153_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N24153_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N24153_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N24153_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C9_N24155_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C9_N24155_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N24155_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N24155_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N24155_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N24155_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N24155_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C17_N24157_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C17_N24157_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N24157_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N24157_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N24157_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N24157_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N24157_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C25_N24159_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C25_N24159_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N24159_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N24159_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N24159_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N24159_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N24159_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C33_N24161_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C33_N24161_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N24161_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N24161_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N24161_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N24161_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N24161_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C41_N24163_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C41_N24163_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N24163_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N24163_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N24163_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N24163_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N24163_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C49_N24165_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C49_N24165_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N24165_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N24165_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N24165_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N24165_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N24165_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C57_N24167_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C57_N24167_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N24167_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N24167_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N24167_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N24167_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N24167_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C65_N24169_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C65_N24169_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N24169_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N24169_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N24169_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N24169_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N24169_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C73_N24171_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C73_N24171_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N24171_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N24171_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N24171_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N24171_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N24171_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [5:0] SBMux_C77_N24215_O_0_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C77_N24215_O_0_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24215_O_0_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24215_O_0_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24215_O_0_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24215_O_0_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N24215_O_0_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C0_N24236_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C0_N24236_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C0_N24236_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C0_N24236_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C0_N24236_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C0_N24236_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C0_N24236_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C8_N24238_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C8_N24238_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C8_N24238_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C8_N24238_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C8_N24238_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C8_N24238_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C8_N24238_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C16_N24240_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C16_N24240_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C16_N24240_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C16_N24240_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C16_N24240_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C16_N24240_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C16_N24240_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C24_N24242_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C24_N24242_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C24_N24242_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C24_N24242_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C24_N24242_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C24_N24242_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C24_N24242_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C32_N24244_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C32_N24244_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C32_N24244_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C32_N24244_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C32_N24244_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C32_N24244_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C32_N24244_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C40_N24246_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C40_N24246_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C40_N24246_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C40_N24246_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C40_N24246_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C40_N24246_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C40_N24246_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C48_N24248_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C48_N24248_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C48_N24248_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C48_N24248_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C48_N24248_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C48_N24248_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C48_N24248_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C56_N24250_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C56_N24250_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C56_N24250_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C56_N24250_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C56_N24250_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C56_N24250_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C56_N24250_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C64_N24252_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C64_N24252_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C64_N24252_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C64_N24252_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C64_N24252_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C64_N24252_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C64_N24252_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C72_N24254_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C72_N24254_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C72_N24254_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C72_N24254_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C72_N24254_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C72_N24254_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C72_N24254_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C76_N24256_O_0_C_4_io_in; // @[TileFull.scala 134:27]
  wire [2:0] SBMux_C76_N24256_O_0_C_4_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N24256_O_0_C_4_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N24256_O_0_C_4_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N24256_O_0_C_4_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N24256_O_0_C_4_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N24256_O_0_C_4_io_arst; // @[TileFull.scala 134:27]
  wire [9:0] SBMux_C1_N28731_O_4_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C1_N28731_O_4_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N28731_O_4_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N28731_O_4_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N28731_O_4_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N28731_O_4_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C1_N28731_O_4_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C9_N28739_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C9_N28739_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N28739_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N28739_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N28739_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N28739_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C9_N28739_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C17_N28747_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C17_N28747_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N28747_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N28747_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N28747_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N28747_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C17_N28747_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C25_N28755_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C25_N28755_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N28755_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N28755_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N28755_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N28755_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C25_N28755_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C33_N28763_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C33_N28763_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N28763_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N28763_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N28763_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N28763_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C33_N28763_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C41_N28771_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C41_N28771_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N28771_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N28771_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N28771_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N28771_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C41_N28771_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C49_N28779_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C49_N28779_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N28779_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N28779_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N28779_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N28779_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C49_N28779_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C57_N28787_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C57_N28787_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N28787_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N28787_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N28787_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N28787_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C57_N28787_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C65_N28795_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C65_N28795_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N28795_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N28795_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N28795_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N28795_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C65_N28795_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C73_N28803_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C73_N28803_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N28803_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N28803_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N28803_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N28803_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C73_N28803_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C77_N28829_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C77_N28829_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N28829_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N28829_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N28829_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N28829_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C77_N28829_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [10:0] SBMux_C0_N28850_O_4_C_7_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C0_N28850_O_4_C_7_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C0_N28850_O_4_C_7_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C0_N28850_O_4_C_7_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C0_N28850_O_4_C_7_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C0_N28850_O_4_C_7_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C0_N28850_O_4_C_7_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C8_N28852_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C8_N28852_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C8_N28852_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C8_N28852_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C8_N28852_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C8_N28852_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C8_N28852_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C16_N28854_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C16_N28854_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C16_N28854_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C16_N28854_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C16_N28854_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C16_N28854_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C16_N28854_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C24_N28856_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C24_N28856_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C24_N28856_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C24_N28856_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C24_N28856_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C24_N28856_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C24_N28856_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C32_N28858_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C32_N28858_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C32_N28858_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C32_N28858_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C32_N28858_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C32_N28858_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C32_N28858_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C40_N28860_O_4_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C40_N28860_O_4_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C40_N28860_O_4_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C40_N28860_O_4_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C40_N28860_O_4_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C40_N28860_O_4_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C40_N28860_O_4_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C48_N28862_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C48_N28862_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C48_N28862_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C48_N28862_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C48_N28862_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C48_N28862_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C48_N28862_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C56_N28864_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C56_N28864_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C56_N28864_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C56_N28864_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C56_N28864_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C56_N28864_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C56_N28864_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [7:0] SBMux_C64_N28866_O_3_C_5_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C64_N28866_O_3_C_5_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C64_N28866_O_3_C_5_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C64_N28866_O_3_C_5_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C64_N28866_O_3_C_5_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C64_N28866_O_3_C_5_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C64_N28866_O_3_C_5_io_arst; // @[TileFull.scala 134:27]
  wire [8:0] SBMux_C72_N28868_O_3_C_6_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C72_N28868_O_3_C_6_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C72_N28868_O_3_C_6_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C72_N28868_O_3_C_6_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C72_N28868_O_3_C_6_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C72_N28868_O_3_C_6_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C72_N28868_O_3_C_6_io_arst; // @[TileFull.scala 134:27]
  wire [9:0] SBMux_C76_N28870_O_3_C_7_io_in; // @[TileFull.scala 134:27]
  wire [3:0] SBMux_C76_N28870_O_3_C_7_io_config; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N28870_O_3_C_7_io_out; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N28870_O_3_C_7_io_loopBreak; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N28870_O_3_C_7_io_ioGndBle; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N28870_O_3_C_7_io_cnstClk; // @[TileFull.scala 134:27]
  wire  SBMux_C76_N28870_O_3_C_7_io_arst; // @[TileFull.scala 134:27]
  wire [4:0] CBMux_IPIN0_N19810_io_in_lo = {IN_CHANY_N28814_20,IN_CHANY_N28741_11,IN_CHANY_N28740_10,IN_CHANY_N28733_3,
    IN_CHANY_N28732_2}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN0_N19810_io_in_hi = {IN_CHANY_N28849_79,IN_CHANY_N28848_78,IN_CHANY_N28837_31,IN_CHANY_N28836_30,
    IN_CHANY_N28815_21}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN1_N19811_io_in_WIRE_1 = SBMux_C25_N28755_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [5:0] CBMux_IPIN1_N19811_io_in_lo = {IN_CHANY_N28813_13,IN_CHANY_N28812_12,IN_CHANY_N28811_5,IN_CHANY_N28810_4,
    _CBMux_IPIN1_N19811_io_in_WIRE_1,IN_CHANY_N28754_24}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN1_N19811_io_in_WIRE_7 = SBMux_C77_N28829_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [5:0] CBMux_IPIN1_N19811_io_in_hi = {IN_CHANY_N28845_63,IN_CHANY_N28844_62,IN_CHANY_N28835_23,IN_CHANY_N28834_22,
    _CBMux_IPIN1_N19811_io_in_WIRE_7,IN_CHANY_N28828_76}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN2_N19812_io_in_WIRE_1 = SBMux_C17_N28747_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [5:0] CBMux_IPIN2_N19812_io_in_lo = {_CBMux_IPIN1_N19811_io_in_WIRE_7,IN_CHANY_N28828_76,IN_CHANY_N28765_35,
    IN_CHANY_N28764_34,_CBMux_IPIN2_N19812_io_in_WIRE_1,IN_CHANY_N28746_16}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN2_N19812_io_in_hi = {IN_CHANY_N28843_55,IN_CHANY_N28842_54,IN_CHANY_N28833_15,IN_CHANY_N28832_14,
    IN_CHANY_N28831_7,IN_CHANY_N28830_6}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN3_N19813_io_in_WIRE_1 = SBMux_C1_N28731_O_4_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN3_N19813_io_in_WIRE_3 = SBMux_C9_N28739_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire [6:0] CBMux_IPIN3_N19813_io_in_lo = {IN_CHANY_N28818_36,IN_CHANY_N28757_27,IN_CHANY_N28756_26,
    _CBMux_IPIN3_N19813_io_in_WIRE_3,IN_CHANY_N28738_8,_CBMux_IPIN3_N19813_io_in_WIRE_1,IN_CHANY_N28730_0}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN3_N19813_io_in_hi = {IN_CHANY_N28849_79,IN_CHANY_N28848_78,IN_CHANY_N28841_47,IN_CHANY_N28840_46,
    IN_CHANY_N28839_39,IN_CHANY_N28838_38,IN_CHANY_N28819_37}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN4_N19814_io_in_WIRE_5 = SBMux_C33_N28763_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [6:0] CBMux_IPIN4_N19814_io_in_lo = {IN_CHANY_N28816_28,_CBMux_IPIN4_N19814_io_in_WIRE_5,IN_CHANY_N28762_32,
    IN_CHANY_N28749_19,IN_CHANY_N28748_18,_CBMux_IPIN3_N19813_io_in_WIRE_1,IN_CHANY_N28730_0}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN4_N19814_io_in_hi = {IN_CHANY_N28849_79,IN_CHANY_N28848_78,IN_CHANY_N28847_71,IN_CHANY_N28846_70,
    IN_CHANY_N28839_39,IN_CHANY_N28838_38,IN_CHANY_N28817_29}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN5_N19815_io_in_lo = {_CBMux_IPIN4_N19814_io_in_WIRE_5,IN_CHANY_N28762_32,IN_CHANY_N28749_19,
    IN_CHANY_N28748_18,IN_CHANY_N28741_11,IN_CHANY_N28740_10}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN5_N19815_io_in_hi = {IN_CHANY_N28847_71,IN_CHANY_N28846_70,_CBMux_IPIN1_N19811_io_in_WIRE_7,
    IN_CHANY_N28828_76,IN_CHANY_N28817_29,IN_CHANY_N28816_28}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN6_N19816_io_in_lo = {IN_CHANY_N28814_20,IN_CHANY_N28813_13,IN_CHANY_N28812_12,IN_CHANY_N28733_3,
    IN_CHANY_N28732_2}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN6_N19816_io_in_hi = {IN_CHANY_N28837_31,IN_CHANY_N28836_30,_CBMux_IPIN1_N19811_io_in_WIRE_7,
    IN_CHANY_N28828_76,IN_CHANY_N28815_21}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN7_N19817_io_in_lo = {IN_CHANY_N28833_15,IN_CHANY_N28832_14,IN_CHANY_N28811_5,IN_CHANY_N28810_4,
    _CBMux_IPIN1_N19811_io_in_WIRE_1,IN_CHANY_N28754_24}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN7_N19817_io_in_hi = {IN_CHANY_N28849_79,IN_CHANY_N28848_78,IN_CHANY_N28845_63,IN_CHANY_N28844_62,
    IN_CHANY_N28835_23,IN_CHANY_N28834_22}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN8_N19818_io_in_lo = {IN_CHANY_N28830_6,IN_CHANY_N28765_35,IN_CHANY_N28764_34,
    _CBMux_IPIN2_N19812_io_in_WIRE_1,IN_CHANY_N28746_16,_CBMux_IPIN3_N19813_io_in_WIRE_3,IN_CHANY_N28738_8}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN8_N19818_io_in_hi = {IN_CHANY_N28849_79,IN_CHANY_N28848_78,IN_CHANY_N28843_55,IN_CHANY_N28842_54,
    IN_CHANY_N28841_47,IN_CHANY_N28840_46,IN_CHANY_N28831_7}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN9_N19819_io_in_lo = {IN_CHANY_N28819_37,IN_CHANY_N28818_36,IN_CHANY_N28757_27,IN_CHANY_N28756_26,
    _CBMux_IPIN3_N19813_io_in_WIRE_3,IN_CHANY_N28738_8}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN9_N19819_io_in_hi = {IN_CHANY_N28841_47,IN_CHANY_N28840_46,IN_CHANY_N28831_7,IN_CHANY_N28830_6,
    _CBMux_IPIN1_N19811_io_in_WIRE_7,IN_CHANY_N28828_76}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN10_N19820_io_in_lo = {IN_CHANY_N28757_27,IN_CHANY_N28756_26,IN_CHANY_N28749_19,IN_CHANY_N28748_18
    ,_CBMux_IPIN3_N19813_io_in_WIRE_1,IN_CHANY_N28730_0}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN10_N19820_io_in_hi = {IN_CHANY_N28839_39,IN_CHANY_N28838_38,_CBMux_IPIN1_N19811_io_in_WIRE_7,
    IN_CHANY_N28828_76,IN_CHANY_N28819_37,IN_CHANY_N28818_36}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN11_N19821_io_in_lo = {IN_CHANY_N28815_21,IN_CHANY_N28814_20,_CBMux_IPIN4_N19814_io_in_WIRE_5,
    IN_CHANY_N28762_32,IN_CHANY_N28741_11,IN_CHANY_N28740_10}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN11_N19821_io_in_hi = {IN_CHANY_N28849_79,IN_CHANY_N28848_78,IN_CHANY_N28847_71,IN_CHANY_N28846_70
    ,IN_CHANY_N28817_29,IN_CHANY_N28816_28}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN12_N19822_io_in_lo = {IN_CHANY_N28834_22,IN_CHANY_N28813_13,IN_CHANY_N28812_12,IN_CHANY_N28733_3,
    IN_CHANY_N28732_2}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN12_N19822_io_in_hi = {IN_CHANY_N28849_79,IN_CHANY_N28848_78,IN_CHANY_N28837_31,IN_CHANY_N28836_30
    ,IN_CHANY_N28835_23}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN13_N19823_io_in_lo = {IN_CHANY_N28828_76,IN_CHANY_N28811_5,IN_CHANY_N28810_4,
    _CBMux_IPIN1_N19811_io_in_WIRE_1,IN_CHANY_N28754_24,_CBMux_IPIN2_N19812_io_in_WIRE_1,IN_CHANY_N28746_16}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN13_N19823_io_in_hi = {IN_CHANY_N28845_63,IN_CHANY_N28844_62,IN_CHANY_N28843_55,IN_CHANY_N28842_54
    ,IN_CHANY_N28833_15,IN_CHANY_N28832_14,_CBMux_IPIN1_N19811_io_in_WIRE_7}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN14_N19824_io_in_lo = {IN_CHANY_N28811_5,IN_CHANY_N28810_4,IN_CHANY_N28765_35,IN_CHANY_N28764_34,
    _CBMux_IPIN2_N19812_io_in_WIRE_1,IN_CHANY_N28746_16}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN14_N19824_io_in_hi = {IN_CHANY_N28843_55,IN_CHANY_N28842_54,IN_CHANY_N28833_15,IN_CHANY_N28832_14
    ,_CBMux_IPIN1_N19811_io_in_WIRE_7,IN_CHANY_N28828_76}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN15_N19825_io_in_lo = {IN_CHANY_N28765_35,IN_CHANY_N28764_34,IN_CHANY_N28757_27,IN_CHANY_N28756_26
    ,_CBMux_IPIN3_N19813_io_in_WIRE_3,IN_CHANY_N28738_8}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN15_N19825_io_in_hi = {IN_CHANY_N28849_79,IN_CHANY_N28848_78,IN_CHANY_N28841_47,IN_CHANY_N28840_46
    ,IN_CHANY_N28831_7,IN_CHANY_N28830_6}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN16_N19826_io_in_WIRE_1 = SBMux_C41_N24163_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN16_N19826_io_in_WIRE_3 = SBMux_C49_N24165_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [5:0] CBMux_IPIN16_N19826_io_in_lo = {IN_CHANX_N24175_3,IN_CHANX_N24174_2,_CBMux_IPIN16_N19826_io_in_WIRE_3,
    IN_CHANX_N24164_48,_CBMux_IPIN16_N19826_io_in_WIRE_1,IN_CHANX_N24162_40}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN16_N19826_io_in_hi = {IN_CHANX_N24223_31,IN_CHANX_N24222_30,IN_CHANX_N24201_21,IN_CHANX_N24200_20
    ,IN_CHANX_N24177_11,IN_CHANX_N24176_10}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN17_N19827_io_in_WIRE_1 = SBMux_C25_N24159_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire [4:0] CBMux_IPIN17_N19827_io_in_lo = {IN_CHANX_N24198_12,IN_CHANX_N24197_5,IN_CHANX_N24196_4,
    _CBMux_IPIN17_N19827_io_in_WIRE_1,IN_CHANX_N24158_24}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN17_N19827_io_in_hi = {IN_CHANX_N24231_63,IN_CHANX_N24230_62,IN_CHANX_N24221_23,IN_CHANX_N24220_22
    ,IN_CHANX_N24199_13}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN18_N19828_io_in_WIRE_1 = SBMux_C17_N24157_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN18_N19828_io_in_WIRE_3 = SBMux_C73_N24171_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire [5:0] CBMux_IPIN18_N19828_io_in_lo = {IN_CHANX_N24183_35,IN_CHANX_N24182_34,_CBMux_IPIN18_N19828_io_in_WIRE_3,
    IN_CHANX_N24170_72,_CBMux_IPIN18_N19828_io_in_WIRE_1,IN_CHANX_N24156_16}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN18_N19828_io_in_hi = {IN_CHANX_N24229_55,IN_CHANX_N24228_54,IN_CHANX_N24219_15,IN_CHANX_N24218_14
    ,IN_CHANX_N24217_7,IN_CHANX_N24216_6}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN19_N19829_io_in_WIRE_1 = SBMux_C1_N24153_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN19_N19829_io_in_WIRE_3 = SBMux_C9_N24155_O_3_C_6_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN19_N19829_io_in_WIRE_5 = SBMux_C65_N24169_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [6:0] CBMux_IPIN19_N19829_io_in_lo = {IN_CHANX_N24180_26,_CBMux_IPIN19_N19829_io_in_WIRE_5,IN_CHANX_N24168_64,
    _CBMux_IPIN19_N19829_io_in_WIRE_3,IN_CHANX_N24154_8,_CBMux_IPIN19_N19829_io_in_WIRE_1,IN_CHANX_N24152_0}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN19_N19829_io_in_hi = {IN_CHANX_N24227_47,IN_CHANX_N24226_46,IN_CHANX_N24225_39,IN_CHANX_N24224_38
    ,IN_CHANX_N24205_37,IN_CHANX_N24204_36,IN_CHANX_N24181_27}; // @[TileFull.scala 166:8]
  wire  _CBMux_IPIN20_N19830_io_in_WIRE_3 = SBMux_C33_N24161_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire  _CBMux_IPIN20_N19830_io_in_WIRE_5 = SBMux_C57_N24167_O_3_C_5_io_out; // @[TileFull.scala 161:{37,37}]
  wire [6:0] CBMux_IPIN20_N19830_io_in_lo = {IN_CHANX_N24178_18,_CBMux_IPIN20_N19830_io_in_WIRE_5,IN_CHANX_N24166_56,
    _CBMux_IPIN20_N19830_io_in_WIRE_3,IN_CHANX_N24160_32,_CBMux_IPIN19_N19829_io_in_WIRE_1,IN_CHANX_N24152_0}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN20_N19830_io_in_hi = {IN_CHANX_N24233_71,IN_CHANX_N24232_70,IN_CHANX_N24225_39,IN_CHANX_N24224_38
    ,IN_CHANX_N24203_29,IN_CHANX_N24202_28,IN_CHANX_N24179_19}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN21_N19831_io_in_lo = {IN_CHANX_N24176_10,_CBMux_IPIN20_N19830_io_in_WIRE_5,IN_CHANX_N24166_56,
    _CBMux_IPIN16_N19826_io_in_WIRE_3,IN_CHANX_N24164_48,_CBMux_IPIN20_N19830_io_in_WIRE_3,IN_CHANX_N24160_32}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN21_N19831_io_in_hi = {IN_CHANX_N24233_71,IN_CHANX_N24232_70,IN_CHANX_N24203_29,IN_CHANX_N24202_28
    ,IN_CHANX_N24179_19,IN_CHANX_N24178_18,IN_CHANX_N24177_11}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN22_N19832_io_in_lo = {IN_CHANX_N24198_12,IN_CHANX_N24175_3,IN_CHANX_N24174_2,
    _CBMux_IPIN16_N19826_io_in_WIRE_1,IN_CHANX_N24162_40}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN22_N19832_io_in_hi = {IN_CHANX_N24223_31,IN_CHANX_N24222_30,IN_CHANX_N24201_21,IN_CHANX_N24200_20
    ,IN_CHANX_N24199_13}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN23_N19833_io_in_lo = {IN_CHANX_N24218_14,IN_CHANX_N24197_5,IN_CHANX_N24196_4,
    _CBMux_IPIN17_N19827_io_in_WIRE_1,IN_CHANX_N24158_24}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN23_N19833_io_in_hi = {IN_CHANX_N24231_63,IN_CHANX_N24230_62,IN_CHANX_N24221_23,IN_CHANX_N24220_22
    ,IN_CHANX_N24219_15}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN24_N19834_io_in_lo = {IN_CHANX_N24182_34,_CBMux_IPIN18_N19828_io_in_WIRE_3,IN_CHANX_N24170_72,
    _CBMux_IPIN18_N19828_io_in_WIRE_1,IN_CHANX_N24156_16,_CBMux_IPIN19_N19829_io_in_WIRE_3,IN_CHANX_N24154_8}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN24_N19834_io_in_hi = {IN_CHANX_N24229_55,IN_CHANX_N24228_54,IN_CHANX_N24227_47,IN_CHANX_N24226_46
    ,IN_CHANX_N24217_7,IN_CHANX_N24216_6,IN_CHANX_N24183_35}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN25_N19835_io_in_lo = {IN_CHANX_N24181_27,IN_CHANX_N24180_26,_CBMux_IPIN19_N19829_io_in_WIRE_5,
    IN_CHANX_N24168_64,_CBMux_IPIN19_N19829_io_in_WIRE_3,IN_CHANX_N24154_8}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN25_N19835_io_in_hi = {IN_CHANX_N24227_47,IN_CHANX_N24226_46,IN_CHANX_N24217_7,IN_CHANX_N24216_6,
    IN_CHANX_N24205_37,IN_CHANX_N24204_36}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN26_N19836_io_in_lo = {IN_CHANX_N24178_18,_CBMux_IPIN19_N19829_io_in_WIRE_5,IN_CHANX_N24168_64,
    _CBMux_IPIN20_N19830_io_in_WIRE_5,IN_CHANX_N24166_56,_CBMux_IPIN19_N19829_io_in_WIRE_1,IN_CHANX_N24152_0}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN26_N19836_io_in_hi = {IN_CHANX_N24225_39,IN_CHANX_N24224_38,IN_CHANX_N24205_37,IN_CHANX_N24204_36
    ,IN_CHANX_N24181_27,IN_CHANX_N24180_26,IN_CHANX_N24179_19}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN27_N19837_io_in_lo = {IN_CHANX_N24177_11,IN_CHANX_N24176_10,_CBMux_IPIN16_N19826_io_in_WIRE_3,
    IN_CHANX_N24164_48,_CBMux_IPIN20_N19830_io_in_WIRE_3,IN_CHANX_N24160_32}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN27_N19837_io_in_hi = {IN_CHANX_N24233_71,IN_CHANX_N24232_70,IN_CHANX_N24203_29,IN_CHANX_N24202_28
    ,IN_CHANX_N24201_21,IN_CHANX_N24200_20}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN28_N19838_io_in_hi = {IN_CHANX_N24223_31,IN_CHANX_N24222_30,IN_CHANX_N24221_23,IN_CHANX_N24220_22
    ,IN_CHANX_N24199_13}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN29_N19839_io_in_lo = {IN_CHANX_N24197_5,IN_CHANX_N24196_4,_CBMux_IPIN17_N19827_io_in_WIRE_1,
    IN_CHANX_N24158_24,_CBMux_IPIN18_N19828_io_in_WIRE_1,IN_CHANX_N24156_16}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN29_N19839_io_in_hi = {IN_CHANX_N24231_63,IN_CHANX_N24230_62,IN_CHANX_N24229_55,IN_CHANX_N24228_54
    ,IN_CHANX_N24219_15,IN_CHANX_N24218_14}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN30_N19840_io_in_hi = {IN_CHANX_N24229_55,IN_CHANX_N24228_54,IN_CHANX_N24219_15,IN_CHANX_N24218_14
    ,IN_CHANX_N24197_5,IN_CHANX_N24196_4}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN31_N19841_io_in_lo = {IN_CHANX_N24180_26,_CBMux_IPIN18_N19828_io_in_WIRE_3,IN_CHANX_N24170_72,
    _CBMux_IPIN19_N19829_io_in_WIRE_5,IN_CHANX_N24168_64,_CBMux_IPIN19_N19829_io_in_WIRE_3,IN_CHANX_N24154_8}; // @[TileFull.scala 166:8]
  wire [6:0] CBMux_IPIN31_N19841_io_in_hi = {IN_CHANX_N24227_47,IN_CHANX_N24226_46,IN_CHANX_N24217_7,IN_CHANX_N24216_6,
    IN_CHANX_N24183_35,IN_CHANX_N24182_34,IN_CHANX_N24181_27}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN32_N19842_io_in_lo = {IN_CHANX_N24179_19,IN_CHANX_N24178_18,_CBMux_IPIN20_N19830_io_in_WIRE_5,
    IN_CHANX_N24166_56,_CBMux_IPIN19_N19829_io_in_WIRE_1,IN_CHANX_N24152_0}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN32_N19842_io_in_hi = {IN_CHANX_N24225_39,IN_CHANX_N24224_38,IN_CHANX_N24205_37,IN_CHANX_N24204_36
    ,IN_CHANX_N24203_29,IN_CHANX_N24202_28}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN33_N19843_io_in_lo = {IN_CHANX_N24176_10,_CBMux_IPIN16_N19826_io_in_WIRE_3,IN_CHANX_N24164_48,
    _CBMux_IPIN20_N19830_io_in_WIRE_3,IN_CHANX_N24160_32}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN33_N19843_io_in_hi = {IN_CHANX_N24223_31,IN_CHANX_N24222_30,IN_CHANX_N24201_21,IN_CHANX_N24200_20
    ,IN_CHANX_N24177_11}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN34_N19844_io_in_lo = {IN_CHANX_N24174_2,_CBMux_IPIN16_N19826_io_in_WIRE_1,IN_CHANX_N24162_40,
    _CBMux_IPIN17_N19827_io_in_WIRE_1,IN_CHANX_N24158_24}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN34_N19844_io_in_hi = {IN_CHANX_N24221_23,IN_CHANX_N24220_22,IN_CHANX_N24199_13,IN_CHANX_N24198_12
    ,IN_CHANX_N24175_3}; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN36_N19846_io_in_lo = {IN_CHANX_N24183_35,IN_CHANX_N24182_34,_CBMux_IPIN18_N19828_io_in_WIRE_1,
    IN_CHANX_N24156_16}; // @[TileFull.scala 166:8]
  wire [3:0] CBMux_IPIN36_N19846_io_in_hi = {IN_CHANX_N24219_15,IN_CHANX_N24218_14,IN_CHANX_N24197_5,IN_CHANX_N24196_4}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN37_N19847_io_in_lo = {IN_CHANX_N24204_36,IN_CHANX_N24181_27,IN_CHANX_N24180_26,
    _CBMux_IPIN19_N19829_io_in_WIRE_3,IN_CHANX_N24154_8}; // @[TileFull.scala 166:8]
  wire [4:0] CBMux_IPIN37_N19847_io_in_hi = {IN_CHANX_N24227_47,IN_CHANX_N24226_46,IN_CHANX_N24217_7,IN_CHANX_N24216_6,
    IN_CHANX_N24205_37}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN38_N19848_io_in_lo = {_CBMux_IPIN20_N19830_io_in_WIRE_5,IN_CHANX_N24166_56,
    _CBMux_IPIN20_N19830_io_in_WIRE_3,IN_CHANX_N24160_32,_CBMux_IPIN19_N19829_io_in_WIRE_1,IN_CHANX_N24152_0}; // @[TileFull.scala 166:8]
  wire [5:0] CBMux_IPIN38_N19848_io_in_hi = {IN_CHANX_N24225_39,IN_CHANX_N24224_38,IN_CHANX_N24203_29,IN_CHANX_N24202_28
    ,IN_CHANX_N24179_19,IN_CHANX_N24178_18}; // @[TileFull.scala 166:8]
  wire  _SBMux_C1_N24153_O_3_C_6_io_in_WIRE_1 = logicBlock_OPIN_51; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C1_N24153_O_3_C_6_io_in_WIRE_0 = logicBlock_OPIN_49; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C1_N24153_O_3_C_6_io_in_WIRE_2 = logicBlock_OPIN_54; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C1_N24153_O_3_C_6_io_in_lo = {IN_CHANX_N24237_1,_SBMux_C1_N24153_O_3_C_6_io_in_WIRE_2,
    _SBMux_C1_N24153_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N24153_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C1_N24153_O_3_C_6_io_in_hi = {IN_CHANY_N28851_1,IN_CHANY_N28837_31,IN_CHANY_N28828_76,
    IN_CHANY_N28816_28,IN_CHANY_N28733_3}; // @[TileFull.scala 183:11]
  wire  _SBMux_C9_N24155_O_3_C_6_io_in_WIRE_1 = logicBlock_OPIN_52; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C9_N24155_O_3_C_6_io_in_lo = {IN_CHANX_N24239_9,_SBMux_C1_N24153_O_3_C_6_io_in_WIRE_2,
    _SBMux_C9_N24155_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N24153_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C9_N24155_O_3_C_6_io_in_hi = {IN_CHANY_N28871_77,IN_CHANY_N28836_30,IN_CHANY_N28817_29,
    IN_CHANY_N28732_2,IN_CHANY_N28730_0}; // @[TileFull.scala 183:11]
  wire  _SBMux_C17_N24157_O_3_C_6_io_in_WIRE_0 = logicBlock_OPIN_50; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C17_N24157_O_3_C_6_io_in_WIRE_2 = logicBlock_OPIN_55; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C17_N24157_O_3_C_6_io_in_lo = {IN_CHANX_N24241_17,_SBMux_C17_N24157_O_3_C_6_io_in_WIRE_2,
    _SBMux_C9_N24155_O_3_C_6_io_in_WIRE_1,_SBMux_C17_N24157_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C17_N24157_O_3_C_6_io_in_hi = {IN_CHANY_N28869_73,IN_CHANY_N28810_4,IN_CHANY_N28764_34,
    IN_CHANY_N28757_27,IN_CHANY_N28738_8}; // @[TileFull.scala 183:11]
  wire  _SBMux_C25_N24159_O_3_C_6_io_in_WIRE_1 = logicBlock_OPIN_53; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C25_N24159_O_3_C_6_io_in_lo = {IN_CHANX_N24243_25,_SBMux_C17_N24157_O_3_C_6_io_in_WIRE_2,
    _SBMux_C25_N24159_O_3_C_6_io_in_WIRE_1,_SBMux_C17_N24157_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C25_N24159_O_3_C_6_io_in_hi = {IN_CHANY_N28867_65,IN_CHANY_N28835_23,IN_CHANY_N28830_6,
    IN_CHANY_N28818_36,IN_CHANY_N28746_16}; // @[TileFull.scala 183:11]
  wire  _SBMux_C33_N24161_O_3_C_5_io_in_WIRE_2 = logicBlock_OPIN_56; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C33_N24161_O_3_C_5_io_in_lo = {IN_CHANX_N24245_33,_SBMux_C33_N24161_O_3_C_5_io_in_WIRE_2,
    _SBMux_C25_N24159_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N24153_O_3_C_6_io_in_WIRE_1}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C33_N24161_O_3_C_5_io_in_hi = {IN_CHANY_N28865_57,IN_CHANY_N28815_21,IN_CHANY_N28754_24,
    IN_CHANY_N28740_10}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C41_N24163_O_3_C_5_io_in_lo = {IN_CHANX_N24247_41,_SBMux_C1_N24153_O_3_C_6_io_in_WIRE_2,
    _SBMux_C1_N24153_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N24153_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C41_N24163_O_3_C_5_io_in_hi = {IN_CHANY_N28863_49,IN_CHANY_N28812_12,IN_CHANY_N28762_32,
    IN_CHANY_N28749_19}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C49_N24165_O_3_C_5_io_in_lo = {IN_CHANX_N24249_49,_SBMux_C1_N24153_O_3_C_6_io_in_WIRE_2,
    _SBMux_C9_N24155_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N24153_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C49_N24165_O_3_C_5_io_in_hi = {IN_CHANY_N28861_41,IN_CHANY_N28833_15,IN_CHANY_N28832_14,
    IN_CHANY_N28770_40}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C57_N24167_O_3_C_5_io_in_lo = {IN_CHANX_N24251_57,_SBMux_C17_N24157_O_3_C_6_io_in_WIRE_2,
    _SBMux_C9_N24155_O_3_C_6_io_in_WIRE_1,_SBMux_C17_N24157_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C57_N24167_O_3_C_5_io_in_hi = {IN_CHANY_N28859_33,IN_CHANY_N28813_13,IN_CHANY_N28778_48,
    IN_CHANY_N28748_18}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C65_N24169_O_3_C_5_io_in_lo = {IN_CHANX_N24253_65,_SBMux_C17_N24157_O_3_C_6_io_in_WIRE_2,
    _SBMux_C25_N24159_O_3_C_6_io_in_WIRE_1,_SBMux_C17_N24157_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C65_N24169_O_3_C_5_io_in_hi = {IN_CHANY_N28857_25,IN_CHANY_N28814_20,IN_CHANY_N28786_56,
    IN_CHANY_N28741_11}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C73_N24171_O_3_C_6_io_in_lo = {IN_CHANX_N24255_73,_SBMux_C33_N24161_O_3_C_5_io_in_WIRE_2,
    _SBMux_C25_N24159_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N24153_O_3_C_6_io_in_WIRE_1}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C73_N24171_O_3_C_6_io_in_hi = {IN_CHANY_N28855_17,IN_CHANY_N28834_22,IN_CHANY_N28831_7,
    IN_CHANY_N28819_37,IN_CHANY_N28794_64}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C77_N24215_O_0_C_6_io_in_lo = {IN_CHANY_N28765_35,IN_CHANY_N28756_26,IN_CHANX_N24257_77}; // @[TileFull.scala 183:11]
  wire [2:0] SBMux_C77_N24215_O_0_C_6_io_in_hi = {IN_CHANY_N28853_9,IN_CHANY_N28811_5,IN_CHANY_N28802_72}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C0_N24236_O_3_C_5_io_in_lo = {IN_CHANX_N24152_0,IN_OPIN_N21024_54,IN_OPIN_N21021_51,IN_OPIN_N21019_49
    }; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C0_N24236_O_3_C_5_io_in_hi = {IN_CHANY_N28871_77,IN_CHANY_N28817_29,IN_CHANY_N28802_72,
    IN_CHANY_N28756_26}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C8_N24238_O_3_C_6_io_in_lo = {IN_CHANX_N24154_8,IN_OPIN_N21024_54,IN_OPIN_N21022_52,IN_OPIN_N21019_49
    }; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C8_N24238_O_3_C_6_io_in_hi = {IN_CHANY_N28851_1,IN_CHANY_N28837_31,IN_CHANY_N28834_22,
    IN_CHANY_N28794_64,IN_CHANY_N28733_3}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C16_N24240_O_3_C_6_io_in_lo = {IN_CHANX_N24156_16,IN_OPIN_N21025_55,IN_OPIN_N21022_52,
    IN_OPIN_N21020_50}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C16_N24240_O_3_C_6_io_in_hi = {IN_CHANY_N28853_9,IN_CHANY_N28814_20,IN_CHANY_N28811_5,
    IN_CHANY_N28786_56,IN_CHANY_N28765_35}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C24_N24242_O_3_C_6_io_in_lo = {IN_CHANX_N24158_24,IN_OPIN_N21025_55,IN_OPIN_N21023_53,
    IN_OPIN_N21020_50}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C24_N24242_O_3_C_6_io_in_hi = {IN_CHANY_N28855_17,IN_CHANY_N28831_7,IN_CHANY_N28819_37,
    IN_CHANY_N28778_48,IN_CHANY_N28748_18}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C32_N24244_O_3_C_5_io_in_lo = {IN_CHANX_N24160_32,IN_OPIN_N21026_56,IN_OPIN_N21023_53,
    IN_OPIN_N21021_51}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C32_N24244_O_3_C_5_io_in_hi = {IN_CHANY_N28857_25,IN_CHANY_N28832_14,IN_CHANY_N28770_40,
    IN_CHANY_N28741_11}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C40_N24246_O_3_C_5_io_in_lo = {IN_CHANX_N24162_40,IN_OPIN_N21024_54,IN_OPIN_N21021_51,
    IN_OPIN_N21019_49}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C40_N24246_O_3_C_5_io_in_hi = {IN_CHANY_N28859_33,IN_CHANY_N28813_13,IN_CHANY_N28812_12,
    IN_CHANY_N28762_32}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C48_N24248_O_3_C_5_io_in_lo = {IN_CHANX_N24164_48,IN_OPIN_N21024_54,IN_OPIN_N21022_52,
    IN_OPIN_N21019_49}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C48_N24248_O_3_C_5_io_in_hi = {IN_CHANY_N28861_41,IN_CHANY_N28833_15,IN_CHANY_N28754_24,
    IN_CHANY_N28740_10}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C56_N24250_O_3_C_5_io_in_lo = {IN_CHANX_N24166_56,IN_OPIN_N21025_55,IN_OPIN_N21022_52,
    IN_OPIN_N21020_50}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C56_N24250_O_3_C_5_io_in_hi = {IN_CHANY_N28863_49,IN_CHANY_N28830_6,IN_CHANY_N28749_19,
    IN_CHANY_N28746_16}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C64_N24252_O_3_C_5_io_in_lo = {IN_CHANX_N24168_64,IN_OPIN_N21025_55,IN_OPIN_N21023_53,
    IN_OPIN_N21020_50}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C64_N24252_O_3_C_5_io_in_hi = {IN_CHANY_N28865_57,IN_CHANY_N28815_21,IN_CHANY_N28810_4,
    IN_CHANY_N28738_8}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C72_N24254_O_3_C_5_io_in_lo = {IN_CHANX_N24170_72,IN_OPIN_N21026_56,IN_OPIN_N21023_53,
    IN_OPIN_N21021_51}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C72_N24254_O_3_C_5_io_in_hi = {IN_CHANY_N28867_65,IN_CHANY_N28835_23,IN_CHANY_N28732_2,
    IN_CHANY_N28730_0}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C76_N24256_O_0_C_4_io_in_lo = {IN_CHANY_N28757_27,IN_CHANX_N24214_76}; // @[TileFull.scala 183:11]
  wire [1:0] SBMux_C76_N24256_O_0_C_4_io_in_hi = {IN_CHANY_N28869_73,IN_CHANY_N28828_76}; // @[TileFull.scala 183:11]
  wire  _SBMux_C1_N28731_O_4_C_6_io_in_WIRE_1 = logicBlock_OPIN_43; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C1_N28731_O_4_C_6_io_in_WIRE_0 = logicBlock_OPIN_41; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C1_N28731_O_4_C_6_io_in_WIRE_3 = logicBlock_OPIN_48; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C1_N28731_O_4_C_6_io_in_WIRE_2 = logicBlock_OPIN_46; // @[TileFull.scala 174:{37,37}]
  wire [4:0] SBMux_C1_N28731_O_4_C_6_io_in_lo = {IN_CHANX_N24154_8,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_3,
    _SBMux_C1_N28731_O_4_C_6_io_in_WIRE_2,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_1,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C1_N28731_O_4_C_6_io_in_hi = {IN_CHANY_N28851_1,IN_CHANX_N24255_73,IN_CHANX_N24196_4,
    IN_CHANX_N24182_34,IN_CHANX_N24181_27}; // @[TileFull.scala 183:11]
  wire  _SBMux_C9_N28739_O_3_C_6_io_in_WIRE_1 = logicBlock_OPIN_44; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C9_N28739_O_3_C_6_io_in_lo = {IN_CHANX_N24156_16,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_2,
    _SBMux_C9_N28739_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C9_N28739_O_3_C_6_io_in_hi = {IN_CHANY_N28853_9,IN_CHANX_N24253_65,IN_CHANX_N24221_23,
    IN_CHANX_N24216_6,IN_CHANX_N24204_36}; // @[TileFull.scala 183:11]
  wire  _SBMux_C17_N28747_O_3_C_5_io_in_WIRE_0 = logicBlock_OPIN_42; // @[TileFull.scala 174:{37,37}]
  wire  _SBMux_C17_N28747_O_3_C_5_io_in_WIRE_2 = logicBlock_OPIN_47; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C17_N28747_O_3_C_5_io_in_lo = {IN_CHANX_N24158_24,_SBMux_C17_N28747_O_3_C_5_io_in_WIRE_2,
    _SBMux_C9_N28739_O_3_C_6_io_in_WIRE_1,_SBMux_C17_N28747_O_3_C_5_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C17_N28747_O_3_C_5_io_in_hi = {IN_CHANY_N28855_17,IN_CHANX_N24251_57,IN_CHANX_N24201_21,
    IN_CHANX_N24176_10}; // @[TileFull.scala 183:11]
  wire  _SBMux_C25_N28755_O_3_C_5_io_in_WIRE_1 = logicBlock_OPIN_45; // @[TileFull.scala 174:{37,37}]
  wire [3:0] SBMux_C25_N28755_O_3_C_5_io_in_lo = {IN_CHANX_N24160_32,_SBMux_C17_N28747_O_3_C_5_io_in_WIRE_2,
    _SBMux_C25_N28755_O_3_C_5_io_in_WIRE_1,_SBMux_C17_N28747_O_3_C_5_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C25_N28755_O_3_C_5_io_in_hi = {IN_CHANY_N28857_25,IN_CHANX_N24249_49,IN_CHANX_N24198_12,
    IN_CHANX_N24179_19}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C33_N28763_O_3_C_5_io_in_lo = {IN_CHANX_N24162_40,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_3,
    _SBMux_C25_N28755_O_3_C_5_io_in_WIRE_1,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_1}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C33_N28763_O_3_C_5_io_in_hi = {IN_CHANY_N28859_33,IN_CHANX_N24247_41,IN_CHANX_N24219_15,
    IN_CHANX_N24218_14}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C41_N28771_O_4_C_5_io_in_lo = {_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_3,
    _SBMux_C1_N28731_O_4_C_6_io_in_WIRE_2,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_1,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C41_N28771_O_4_C_5_io_in_hi = {IN_CHANY_N28861_41,IN_CHANX_N24245_33,IN_CHANX_N24199_13,
    IN_CHANX_N24178_18,IN_CHANX_N24164_48}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C49_N28779_O_3_C_5_io_in_lo = {IN_CHANX_N24166_56,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_2,
    _SBMux_C9_N28739_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C49_N28779_O_3_C_5_io_in_hi = {IN_CHANY_N28863_49,IN_CHANX_N24243_25,IN_CHANX_N24200_20,
    IN_CHANX_N24177_11}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C57_N28787_O_3_C_5_io_in_lo = {IN_CHANX_N24168_64,_SBMux_C17_N28747_O_3_C_5_io_in_WIRE_2,
    _SBMux_C9_N28739_O_3_C_6_io_in_WIRE_1,_SBMux_C17_N28747_O_3_C_5_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C57_N28787_O_3_C_5_io_in_hi = {IN_CHANY_N28865_57,IN_CHANX_N24241_17,IN_CHANX_N24220_22,
    IN_CHANX_N24217_7}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C65_N28795_O_3_C_5_io_in_lo = {IN_CHANX_N24170_72,_SBMux_C17_N28747_O_3_C_5_io_in_WIRE_2,
    _SBMux_C25_N28755_O_3_C_5_io_in_WIRE_1,_SBMux_C17_N28747_O_3_C_5_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C65_N28795_O_3_C_5_io_in_hi = {IN_CHANY_N28867_65,IN_CHANX_N24239_9,IN_CHANX_N24197_5,
    IN_CHANX_N24180_26}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C73_N28803_O_3_C_5_io_in_lo = {IN_CHANX_N24175_3,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_3,
    _SBMux_C25_N28755_O_3_C_5_io_in_WIRE_1,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_1}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C73_N28803_O_3_C_5_io_in_hi = {IN_CHANY_N28869_73,IN_CHANX_N24237_1,IN_CHANX_N24214_76,
    IN_CHANX_N24202_28}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C77_N28829_O_3_C_5_io_in_lo = {IN_CHANX_N24152_0,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_1,
    _SBMux_C17_N28747_O_3_C_5_io_in_WIRE_0,_SBMux_C1_N28731_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C77_N28829_O_3_C_5_io_in_hi = {IN_CHANY_N28871_77,IN_CHANX_N24257_77,IN_CHANX_N24222_30,
    IN_CHANX_N24174_2}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C0_N28850_O_4_C_7_io_in_lo = {IN_CHANX_N24152_0,IN_OPIN_N19974_48,IN_OPIN_N19972_46,IN_OPIN_N19969_43
    ,IN_OPIN_N19967_41}; // @[TileFull.scala 183:11]
  wire [5:0] SBMux_C0_N28850_O_4_C_7_io_in_hi = {IN_CHANY_N28730_0,IN_CHANX_N24239_9,IN_CHANX_N24222_30,
    IN_CHANX_N24197_5,IN_CHANX_N24183_35,IN_CHANX_N24174_2}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C8_N28852_O_3_C_6_io_in_lo = {IN_CHANX_N24202_28,IN_OPIN_N19972_46,IN_OPIN_N19970_44,
    IN_OPIN_N19967_41}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C8_N28852_O_3_C_6_io_in_hi = {IN_CHANY_N28738_8,IN_CHANX_N24241_17,IN_CHANX_N24217_7,
    IN_CHANX_N24214_76,IN_CHANX_N24205_37}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C16_N28854_O_3_C_5_io_in_lo = {IN_CHANX_N24170_72,IN_OPIN_N19973_47,IN_OPIN_N19970_44,
    IN_OPIN_N19968_42}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C16_N28854_O_3_C_5_io_in_hi = {IN_CHANY_N28746_16,IN_CHANX_N24243_25,IN_CHANX_N24180_26,
    IN_CHANX_N24177_11}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C24_N28856_O_3_C_5_io_in_lo = {IN_CHANX_N24168_64,IN_OPIN_N19973_47,IN_OPIN_N19971_45,
    IN_OPIN_N19968_42}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C24_N28856_O_3_C_5_io_in_hi = {IN_CHANY_N28754_24,IN_CHANX_N24245_33,IN_CHANX_N24220_22,
    IN_CHANX_N24199_13}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C32_N28858_O_3_C_5_io_in_lo = {IN_CHANX_N24166_56,IN_OPIN_N19974_48,IN_OPIN_N19971_45,
    IN_OPIN_N19969_43}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C32_N28858_O_3_C_5_io_in_hi = {IN_CHANY_N28762_32,IN_CHANX_N24247_41,IN_CHANX_N24219_15,
    IN_CHANX_N24200_20}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C40_N28860_O_4_C_5_io_in_lo = {IN_OPIN_N19974_48,IN_OPIN_N19972_46,IN_OPIN_N19969_43,
    IN_OPIN_N19967_41}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C40_N28860_O_4_C_5_io_in_hi = {IN_CHANY_N28770_40,IN_CHANX_N24249_49,IN_CHANX_N24179_19,
    IN_CHANX_N24178_18,IN_CHANX_N24164_48}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C48_N28862_O_3_C_5_io_in_lo = {IN_CHANX_N24162_40,IN_OPIN_N19972_46,IN_OPIN_N19970_44,
    IN_OPIN_N19967_41}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C48_N28862_O_3_C_5_io_in_hi = {IN_CHANY_N28778_48,IN_CHANX_N24251_57,IN_CHANX_N24218_14,
    IN_CHANX_N24201_21}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C56_N28864_O_3_C_5_io_in_lo = {IN_CHANX_N24160_32,IN_OPIN_N19973_47,IN_OPIN_N19970_44,
    IN_OPIN_N19968_42}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C56_N28864_O_3_C_5_io_in_hi = {IN_CHANY_N28786_56,IN_CHANX_N24253_65,IN_CHANX_N24221_23,
    IN_CHANX_N24198_12}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C64_N28866_O_3_C_5_io_in_lo = {IN_CHANX_N24158_24,IN_OPIN_N19973_47,IN_OPIN_N19971_45,
    IN_OPIN_N19968_42}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C64_N28866_O_3_C_5_io_in_hi = {IN_CHANY_N28794_64,IN_CHANX_N24255_73,IN_CHANX_N24181_27,
    IN_CHANX_N24176_10}; // @[TileFull.scala 183:11]
  wire [3:0] SBMux_C72_N28868_O_3_C_6_io_in_lo = {IN_CHANX_N24156_16,IN_OPIN_N19974_48,IN_OPIN_N19971_45,
    IN_OPIN_N19969_43}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C72_N28868_O_3_C_6_io_in_hi = {IN_CHANY_N28802_72,IN_CHANX_N24257_77,IN_CHANX_N24216_6,
    IN_CHANX_N24204_36,IN_CHANX_N24203_29}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C76_N28870_O_3_C_7_io_in_lo = {IN_CHANX_N24175_3,IN_CHANX_N24154_8,IN_OPIN_N19969_43,
    IN_OPIN_N19968_42,IN_OPIN_N19967_41}; // @[TileFull.scala 183:11]
  wire [4:0] SBMux_C76_N28870_O_3_C_7_io_in_hi = {IN_CHANY_N28828_76,IN_CHANX_N24237_1,IN_CHANX_N24223_31,
    IN_CHANX_N24196_4,IN_CHANX_N24182_34}; // @[TileFull.scala 183:11]
  CLBlut4N10Mem logicBlock ( // @[TileFull.scala 46:37]
    .IPIN_0(logicBlock_IPIN_0),
    .IPIN_1(logicBlock_IPIN_1),
    .IPIN_2(logicBlock_IPIN_2),
    .IPIN_3(logicBlock_IPIN_3),
    .IPIN_4(logicBlock_IPIN_4),
    .IPIN_5(logicBlock_IPIN_5),
    .IPIN_6(logicBlock_IPIN_6),
    .IPIN_7(logicBlock_IPIN_7),
    .IPIN_8(logicBlock_IPIN_8),
    .IPIN_9(logicBlock_IPIN_9),
    .IPIN_10(logicBlock_IPIN_10),
    .IPIN_11(logicBlock_IPIN_11),
    .IPIN_12(logicBlock_IPIN_12),
    .IPIN_13(logicBlock_IPIN_13),
    .IPIN_14(logicBlock_IPIN_14),
    .IPIN_15(logicBlock_IPIN_15),
    .IPIN_16(logicBlock_IPIN_16),
    .IPIN_17(logicBlock_IPIN_17),
    .IPIN_18(logicBlock_IPIN_18),
    .IPIN_19(logicBlock_IPIN_19),
    .IPIN_20(logicBlock_IPIN_20),
    .IPIN_21(logicBlock_IPIN_21),
    .IPIN_22(logicBlock_IPIN_22),
    .IPIN_23(logicBlock_IPIN_23),
    .IPIN_24(logicBlock_IPIN_24),
    .IPIN_25(logicBlock_IPIN_25),
    .IPIN_26(logicBlock_IPIN_26),
    .IPIN_27(logicBlock_IPIN_27),
    .IPIN_28(logicBlock_IPIN_28),
    .IPIN_29(logicBlock_IPIN_29),
    .IPIN_30(logicBlock_IPIN_30),
    .IPIN_31(logicBlock_IPIN_31),
    .OPIN_41(logicBlock_OPIN_41),
    .OPIN_42(logicBlock_OPIN_42),
    .OPIN_43(logicBlock_OPIN_43),
    .OPIN_44(logicBlock_OPIN_44),
    .OPIN_45(logicBlock_OPIN_45),
    .OPIN_46(logicBlock_OPIN_46),
    .OPIN_47(logicBlock_OPIN_47),
    .OPIN_48(logicBlock_OPIN_48),
    .OPIN_49(logicBlock_OPIN_49),
    .OPIN_50(logicBlock_OPIN_50),
    .OPIN_51(logicBlock_OPIN_51),
    .OPIN_52(logicBlock_OPIN_52),
    .OPIN_53(logicBlock_OPIN_53),
    .OPIN_54(logicBlock_OPIN_54),
    .OPIN_55(logicBlock_OPIN_55),
    .OPIN_56(logicBlock_OPIN_56),
    .clock(logicBlock_clock),
    .reset(logicBlock_reset),
    .ioPad_i(logicBlock_ioPad_i),
    .configBits(logicBlock_configBits),
    .gndLBouts(logicBlock_gndLBouts)
  );
  ScanConf_Tile_9_3_clbmemtile configBlock ( // @[TileFull.scala 61:31]
    .clock(configBlock_clock),
    .ioBundle_confOut(configBlock_ioBundle_confOut),
    .ioBundle_scan_in(configBlock_ioBundle_scan_in),
    .ioBundle_scan_en(configBlock_ioBundle_scan_en),
    .ioBundle_scan_out(configBlock_ioBundle_scan_out)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN0_N19810 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN0_N19810_io_in),
    .io_config(CBMux_IPIN0_N19810_io_config),
    .io_out(CBMux_IPIN0_N19810_io_out),
    .io_loopBreak(CBMux_IPIN0_N19810_io_loopBreak),
    .io_cnstClk(CBMux_IPIN0_N19810_io_cnstClk),
    .io_arst(CBMux_IPIN0_N19810_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN1_N19811 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN1_N19811_io_in),
    .io_config(CBMux_IPIN1_N19811_io_config),
    .io_out(CBMux_IPIN1_N19811_io_out),
    .io_loopBreak(CBMux_IPIN1_N19811_io_loopBreak),
    .io_cnstClk(CBMux_IPIN1_N19811_io_cnstClk),
    .io_arst(CBMux_IPIN1_N19811_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN2_N19812 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN2_N19812_io_in),
    .io_config(CBMux_IPIN2_N19812_io_config),
    .io_out(CBMux_IPIN2_N19812_io_out),
    .io_loopBreak(CBMux_IPIN2_N19812_io_loopBreak),
    .io_cnstClk(CBMux_IPIN2_N19812_io_cnstClk),
    .io_arst(CBMux_IPIN2_N19812_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN3_N19813 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN3_N19813_io_in),
    .io_config(CBMux_IPIN3_N19813_io_config),
    .io_out(CBMux_IPIN3_N19813_io_out),
    .io_loopBreak(CBMux_IPIN3_N19813_io_loopBreak),
    .io_cnstClk(CBMux_IPIN3_N19813_io_cnstClk),
    .io_arst(CBMux_IPIN3_N19813_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN4_N19814 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN4_N19814_io_in),
    .io_config(CBMux_IPIN4_N19814_io_config),
    .io_out(CBMux_IPIN4_N19814_io_out),
    .io_loopBreak(CBMux_IPIN4_N19814_io_loopBreak),
    .io_cnstClk(CBMux_IPIN4_N19814_io_cnstClk),
    .io_arst(CBMux_IPIN4_N19814_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN5_N19815 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN5_N19815_io_in),
    .io_config(CBMux_IPIN5_N19815_io_config),
    .io_out(CBMux_IPIN5_N19815_io_out),
    .io_loopBreak(CBMux_IPIN5_N19815_io_loopBreak),
    .io_cnstClk(CBMux_IPIN5_N19815_io_cnstClk),
    .io_arst(CBMux_IPIN5_N19815_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN6_N19816 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN6_N19816_io_in),
    .io_config(CBMux_IPIN6_N19816_io_config),
    .io_out(CBMux_IPIN6_N19816_io_out),
    .io_loopBreak(CBMux_IPIN6_N19816_io_loopBreak),
    .io_cnstClk(CBMux_IPIN6_N19816_io_cnstClk),
    .io_arst(CBMux_IPIN6_N19816_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN7_N19817 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN7_N19817_io_in),
    .io_config(CBMux_IPIN7_N19817_io_config),
    .io_out(CBMux_IPIN7_N19817_io_out),
    .io_loopBreak(CBMux_IPIN7_N19817_io_loopBreak),
    .io_cnstClk(CBMux_IPIN7_N19817_io_cnstClk),
    .io_arst(CBMux_IPIN7_N19817_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN8_N19818 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN8_N19818_io_in),
    .io_config(CBMux_IPIN8_N19818_io_config),
    .io_out(CBMux_IPIN8_N19818_io_out),
    .io_loopBreak(CBMux_IPIN8_N19818_io_loopBreak),
    .io_cnstClk(CBMux_IPIN8_N19818_io_cnstClk),
    .io_arst(CBMux_IPIN8_N19818_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN9_N19819 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN9_N19819_io_in),
    .io_config(CBMux_IPIN9_N19819_io_config),
    .io_out(CBMux_IPIN9_N19819_io_out),
    .io_loopBreak(CBMux_IPIN9_N19819_io_loopBreak),
    .io_cnstClk(CBMux_IPIN9_N19819_io_cnstClk),
    .io_arst(CBMux_IPIN9_N19819_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN10_N19820 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN10_N19820_io_in),
    .io_config(CBMux_IPIN10_N19820_io_config),
    .io_out(CBMux_IPIN10_N19820_io_out),
    .io_loopBreak(CBMux_IPIN10_N19820_io_loopBreak),
    .io_cnstClk(CBMux_IPIN10_N19820_io_cnstClk),
    .io_arst(CBMux_IPIN10_N19820_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN11_N19821 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN11_N19821_io_in),
    .io_config(CBMux_IPIN11_N19821_io_config),
    .io_out(CBMux_IPIN11_N19821_io_out),
    .io_loopBreak(CBMux_IPIN11_N19821_io_loopBreak),
    .io_cnstClk(CBMux_IPIN11_N19821_io_cnstClk),
    .io_arst(CBMux_IPIN11_N19821_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN12_N19822 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN12_N19822_io_in),
    .io_config(CBMux_IPIN12_N19822_io_config),
    .io_out(CBMux_IPIN12_N19822_io_out),
    .io_loopBreak(CBMux_IPIN12_N19822_io_loopBreak),
    .io_cnstClk(CBMux_IPIN12_N19822_io_cnstClk),
    .io_arst(CBMux_IPIN12_N19822_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN13_N19823 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN13_N19823_io_in),
    .io_config(CBMux_IPIN13_N19823_io_config),
    .io_out(CBMux_IPIN13_N19823_io_out),
    .io_loopBreak(CBMux_IPIN13_N19823_io_loopBreak),
    .io_cnstClk(CBMux_IPIN13_N19823_io_cnstClk),
    .io_arst(CBMux_IPIN13_N19823_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN14_N19824 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN14_N19824_io_in),
    .io_config(CBMux_IPIN14_N19824_io_config),
    .io_out(CBMux_IPIN14_N19824_io_out),
    .io_loopBreak(CBMux_IPIN14_N19824_io_loopBreak),
    .io_cnstClk(CBMux_IPIN14_N19824_io_cnstClk),
    .io_arst(CBMux_IPIN14_N19824_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN15_N19825 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN15_N19825_io_in),
    .io_config(CBMux_IPIN15_N19825_io_config),
    .io_out(CBMux_IPIN15_N19825_io_out),
    .io_loopBreak(CBMux_IPIN15_N19825_io_loopBreak),
    .io_cnstClk(CBMux_IPIN15_N19825_io_cnstClk),
    .io_arst(CBMux_IPIN15_N19825_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN16_N19826 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN16_N19826_io_in),
    .io_config(CBMux_IPIN16_N19826_io_config),
    .io_out(CBMux_IPIN16_N19826_io_out),
    .io_loopBreak(CBMux_IPIN16_N19826_io_loopBreak),
    .io_cnstClk(CBMux_IPIN16_N19826_io_cnstClk),
    .io_arst(CBMux_IPIN16_N19826_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN17_N19827 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN17_N19827_io_in),
    .io_config(CBMux_IPIN17_N19827_io_config),
    .io_out(CBMux_IPIN17_N19827_io_out),
    .io_loopBreak(CBMux_IPIN17_N19827_io_loopBreak),
    .io_cnstClk(CBMux_IPIN17_N19827_io_cnstClk),
    .io_arst(CBMux_IPIN17_N19827_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN18_N19828 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN18_N19828_io_in),
    .io_config(CBMux_IPIN18_N19828_io_config),
    .io_out(CBMux_IPIN18_N19828_io_out),
    .io_loopBreak(CBMux_IPIN18_N19828_io_loopBreak),
    .io_cnstClk(CBMux_IPIN18_N19828_io_cnstClk),
    .io_arst(CBMux_IPIN18_N19828_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN19_N19829 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN19_N19829_io_in),
    .io_config(CBMux_IPIN19_N19829_io_config),
    .io_out(CBMux_IPIN19_N19829_io_out),
    .io_loopBreak(CBMux_IPIN19_N19829_io_loopBreak),
    .io_cnstClk(CBMux_IPIN19_N19829_io_cnstClk),
    .io_arst(CBMux_IPIN19_N19829_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN20_N19830 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN20_N19830_io_in),
    .io_config(CBMux_IPIN20_N19830_io_config),
    .io_out(CBMux_IPIN20_N19830_io_out),
    .io_loopBreak(CBMux_IPIN20_N19830_io_loopBreak),
    .io_cnstClk(CBMux_IPIN20_N19830_io_cnstClk),
    .io_arst(CBMux_IPIN20_N19830_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN21_N19831 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN21_N19831_io_in),
    .io_config(CBMux_IPIN21_N19831_io_config),
    .io_out(CBMux_IPIN21_N19831_io_out),
    .io_loopBreak(CBMux_IPIN21_N19831_io_loopBreak),
    .io_cnstClk(CBMux_IPIN21_N19831_io_cnstClk),
    .io_arst(CBMux_IPIN21_N19831_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN22_N19832 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN22_N19832_io_in),
    .io_config(CBMux_IPIN22_N19832_io_config),
    .io_out(CBMux_IPIN22_N19832_io_out),
    .io_loopBreak(CBMux_IPIN22_N19832_io_loopBreak),
    .io_cnstClk(CBMux_IPIN22_N19832_io_cnstClk),
    .io_arst(CBMux_IPIN22_N19832_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN23_N19833 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN23_N19833_io_in),
    .io_config(CBMux_IPIN23_N19833_io_config),
    .io_out(CBMux_IPIN23_N19833_io_out),
    .io_loopBreak(CBMux_IPIN23_N19833_io_loopBreak),
    .io_cnstClk(CBMux_IPIN23_N19833_io_cnstClk),
    .io_arst(CBMux_IPIN23_N19833_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN24_N19834 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN24_N19834_io_in),
    .io_config(CBMux_IPIN24_N19834_io_config),
    .io_out(CBMux_IPIN24_N19834_io_out),
    .io_loopBreak(CBMux_IPIN24_N19834_io_loopBreak),
    .io_cnstClk(CBMux_IPIN24_N19834_io_cnstClk),
    .io_arst(CBMux_IPIN24_N19834_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN25_N19835 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN25_N19835_io_in),
    .io_config(CBMux_IPIN25_N19835_io_config),
    .io_out(CBMux_IPIN25_N19835_io_out),
    .io_loopBreak(CBMux_IPIN25_N19835_io_loopBreak),
    .io_cnstClk(CBMux_IPIN25_N19835_io_cnstClk),
    .io_arst(CBMux_IPIN25_N19835_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN26_N19836 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN26_N19836_io_in),
    .io_config(CBMux_IPIN26_N19836_io_config),
    .io_out(CBMux_IPIN26_N19836_io_out),
    .io_loopBreak(CBMux_IPIN26_N19836_io_loopBreak),
    .io_cnstClk(CBMux_IPIN26_N19836_io_cnstClk),
    .io_arst(CBMux_IPIN26_N19836_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN27_N19837 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN27_N19837_io_in),
    .io_config(CBMux_IPIN27_N19837_io_config),
    .io_out(CBMux_IPIN27_N19837_io_out),
    .io_loopBreak(CBMux_IPIN27_N19837_io_loopBreak),
    .io_cnstClk(CBMux_IPIN27_N19837_io_cnstClk),
    .io_arst(CBMux_IPIN27_N19837_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN28_N19838 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN28_N19838_io_in),
    .io_config(CBMux_IPIN28_N19838_io_config),
    .io_out(CBMux_IPIN28_N19838_io_out),
    .io_loopBreak(CBMux_IPIN28_N19838_io_loopBreak),
    .io_cnstClk(CBMux_IPIN28_N19838_io_cnstClk),
    .io_arst(CBMux_IPIN28_N19838_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN29_N19839 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN29_N19839_io_in),
    .io_config(CBMux_IPIN29_N19839_io_config),
    .io_out(CBMux_IPIN29_N19839_io_out),
    .io_loopBreak(CBMux_IPIN29_N19839_io_loopBreak),
    .io_cnstClk(CBMux_IPIN29_N19839_io_cnstClk),
    .io_arst(CBMux_IPIN29_N19839_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN30_N19840 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN30_N19840_io_in),
    .io_config(CBMux_IPIN30_N19840_io_config),
    .io_out(CBMux_IPIN30_N19840_io_out),
    .io_loopBreak(CBMux_IPIN30_N19840_io_loopBreak),
    .io_cnstClk(CBMux_IPIN30_N19840_io_cnstClk),
    .io_arst(CBMux_IPIN30_N19840_io_arst)
  );
  MuxNInput_14_SCAOptCB CBMux_IPIN31_N19841 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN31_N19841_io_in),
    .io_config(CBMux_IPIN31_N19841_io_config),
    .io_out(CBMux_IPIN31_N19841_io_out),
    .io_loopBreak(CBMux_IPIN31_N19841_io_loopBreak),
    .io_cnstClk(CBMux_IPIN31_N19841_io_cnstClk),
    .io_arst(CBMux_IPIN31_N19841_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN32_N19842 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN32_N19842_io_in),
    .io_config(CBMux_IPIN32_N19842_io_config),
    .io_out(CBMux_IPIN32_N19842_io_out),
    .io_loopBreak(CBMux_IPIN32_N19842_io_loopBreak),
    .io_cnstClk(CBMux_IPIN32_N19842_io_cnstClk),
    .io_arst(CBMux_IPIN32_N19842_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN33_N19843 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN33_N19843_io_in),
    .io_config(CBMux_IPIN33_N19843_io_config),
    .io_out(CBMux_IPIN33_N19843_io_out),
    .io_loopBreak(CBMux_IPIN33_N19843_io_loopBreak),
    .io_cnstClk(CBMux_IPIN33_N19843_io_cnstClk),
    .io_arst(CBMux_IPIN33_N19843_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN34_N19844 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN34_N19844_io_in),
    .io_config(CBMux_IPIN34_N19844_io_config),
    .io_out(CBMux_IPIN34_N19844_io_out),
    .io_loopBreak(CBMux_IPIN34_N19844_io_loopBreak),
    .io_cnstClk(CBMux_IPIN34_N19844_io_cnstClk),
    .io_arst(CBMux_IPIN34_N19844_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN35_N19845 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN35_N19845_io_in),
    .io_config(CBMux_IPIN35_N19845_io_config),
    .io_out(CBMux_IPIN35_N19845_io_out),
    .io_loopBreak(CBMux_IPIN35_N19845_io_loopBreak),
    .io_cnstClk(CBMux_IPIN35_N19845_io_cnstClk),
    .io_arst(CBMux_IPIN35_N19845_io_arst)
  );
  MuxNInput_8_SCAOptCB CBMux_IPIN36_N19846 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN36_N19846_io_in),
    .io_config(CBMux_IPIN36_N19846_io_config),
    .io_loopBreak(CBMux_IPIN36_N19846_io_loopBreak),
    .io_cnstClk(CBMux_IPIN36_N19846_io_cnstClk),
    .io_arst(CBMux_IPIN36_N19846_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN37_N19847 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN37_N19847_io_in),
    .io_config(CBMux_IPIN37_N19847_io_config),
    .io_out(CBMux_IPIN37_N19847_io_out),
    .io_loopBreak(CBMux_IPIN37_N19847_io_loopBreak),
    .io_cnstClk(CBMux_IPIN37_N19847_io_cnstClk),
    .io_arst(CBMux_IPIN37_N19847_io_arst)
  );
  MuxNInput_12_SCAOptCB CBMux_IPIN38_N19848 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN38_N19848_io_in),
    .io_config(CBMux_IPIN38_N19848_io_config),
    .io_out(CBMux_IPIN38_N19848_io_out),
    .io_loopBreak(CBMux_IPIN38_N19848_io_loopBreak),
    .io_cnstClk(CBMux_IPIN38_N19848_io_cnstClk),
    .io_arst(CBMux_IPIN38_N19848_io_arst)
  );
  MuxNInput_10_SCAOptCB CBMux_IPIN39_N19849 ( // @[TileFull.scala 97:27]
    .io_in(CBMux_IPIN39_N19849_io_in),
    .io_config(CBMux_IPIN39_N19849_io_config),
    .io_out(CBMux_IPIN39_N19849_io_out),
    .io_loopBreak(CBMux_IPIN39_N19849_io_loopBreak),
    .io_cnstClk(CBMux_IPIN39_N19849_io_cnstClk),
    .io_arst(CBMux_IPIN39_N19849_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C1_N24153_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C1_N24153_O_3_C_6_io_in),
    .io_config(SBMux_C1_N24153_O_3_C_6_io_config),
    .io_out(SBMux_C1_N24153_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C1_N24153_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C1_N24153_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C1_N24153_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C1_N24153_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C9_N24155_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C9_N24155_O_3_C_6_io_in),
    .io_config(SBMux_C9_N24155_O_3_C_6_io_config),
    .io_out(SBMux_C9_N24155_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C9_N24155_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C9_N24155_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C9_N24155_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C9_N24155_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C17_N24157_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C17_N24157_O_3_C_6_io_in),
    .io_config(SBMux_C17_N24157_O_3_C_6_io_config),
    .io_out(SBMux_C17_N24157_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C17_N24157_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C17_N24157_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C17_N24157_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C17_N24157_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C25_N24159_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C25_N24159_O_3_C_6_io_in),
    .io_config(SBMux_C25_N24159_O_3_C_6_io_config),
    .io_out(SBMux_C25_N24159_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C25_N24159_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C25_N24159_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C25_N24159_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C25_N24159_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C33_N24161_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C33_N24161_O_3_C_5_io_in),
    .io_config(SBMux_C33_N24161_O_3_C_5_io_config),
    .io_out(SBMux_C33_N24161_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C33_N24161_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C33_N24161_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C33_N24161_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C33_N24161_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C41_N24163_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C41_N24163_O_3_C_5_io_in),
    .io_config(SBMux_C41_N24163_O_3_C_5_io_config),
    .io_out(SBMux_C41_N24163_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C41_N24163_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C41_N24163_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C41_N24163_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C41_N24163_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C49_N24165_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C49_N24165_O_3_C_5_io_in),
    .io_config(SBMux_C49_N24165_O_3_C_5_io_config),
    .io_out(SBMux_C49_N24165_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C49_N24165_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C49_N24165_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C49_N24165_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C49_N24165_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C57_N24167_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C57_N24167_O_3_C_5_io_in),
    .io_config(SBMux_C57_N24167_O_3_C_5_io_config),
    .io_out(SBMux_C57_N24167_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C57_N24167_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C57_N24167_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C57_N24167_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C57_N24167_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C65_N24169_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C65_N24169_O_3_C_5_io_in),
    .io_config(SBMux_C65_N24169_O_3_C_5_io_config),
    .io_out(SBMux_C65_N24169_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C65_N24169_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C65_N24169_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C65_N24169_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C65_N24169_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C73_N24171_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C73_N24171_O_3_C_6_io_in),
    .io_config(SBMux_C73_N24171_O_3_C_6_io_config),
    .io_out(SBMux_C73_N24171_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C73_N24171_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C73_N24171_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C73_N24171_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C73_N24171_O_3_C_6_io_arst)
  );
  MuxNInput_O0_C6_SCAOptSB SBMux_C77_N24215_O_0_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C77_N24215_O_0_C_6_io_in),
    .io_config(SBMux_C77_N24215_O_0_C_6_io_config),
    .io_out(SBMux_C77_N24215_O_0_C_6_io_out),
    .io_loopBreak(SBMux_C77_N24215_O_0_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C77_N24215_O_0_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C77_N24215_O_0_C_6_io_cnstClk),
    .io_arst(SBMux_C77_N24215_O_0_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C0_N24236_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C0_N24236_O_3_C_5_io_in),
    .io_config(SBMux_C0_N24236_O_3_C_5_io_config),
    .io_out(SBMux_C0_N24236_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C0_N24236_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C0_N24236_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C0_N24236_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C0_N24236_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C8_N24238_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C8_N24238_O_3_C_6_io_in),
    .io_config(SBMux_C8_N24238_O_3_C_6_io_config),
    .io_out(SBMux_C8_N24238_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C8_N24238_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C8_N24238_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C8_N24238_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C8_N24238_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C16_N24240_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C16_N24240_O_3_C_6_io_in),
    .io_config(SBMux_C16_N24240_O_3_C_6_io_config),
    .io_out(SBMux_C16_N24240_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C16_N24240_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C16_N24240_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C16_N24240_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C16_N24240_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C24_N24242_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C24_N24242_O_3_C_6_io_in),
    .io_config(SBMux_C24_N24242_O_3_C_6_io_config),
    .io_out(SBMux_C24_N24242_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C24_N24242_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C24_N24242_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C24_N24242_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C24_N24242_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C32_N24244_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C32_N24244_O_3_C_5_io_in),
    .io_config(SBMux_C32_N24244_O_3_C_5_io_config),
    .io_out(SBMux_C32_N24244_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C32_N24244_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C32_N24244_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C32_N24244_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C32_N24244_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C40_N24246_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C40_N24246_O_3_C_5_io_in),
    .io_config(SBMux_C40_N24246_O_3_C_5_io_config),
    .io_out(SBMux_C40_N24246_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C40_N24246_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C40_N24246_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C40_N24246_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C40_N24246_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C48_N24248_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C48_N24248_O_3_C_5_io_in),
    .io_config(SBMux_C48_N24248_O_3_C_5_io_config),
    .io_out(SBMux_C48_N24248_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C48_N24248_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C48_N24248_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C48_N24248_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C48_N24248_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C56_N24250_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C56_N24250_O_3_C_5_io_in),
    .io_config(SBMux_C56_N24250_O_3_C_5_io_config),
    .io_out(SBMux_C56_N24250_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C56_N24250_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C56_N24250_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C56_N24250_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C56_N24250_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C64_N24252_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C64_N24252_O_3_C_5_io_in),
    .io_config(SBMux_C64_N24252_O_3_C_5_io_config),
    .io_out(SBMux_C64_N24252_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C64_N24252_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C64_N24252_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C64_N24252_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C64_N24252_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C72_N24254_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C72_N24254_O_3_C_5_io_in),
    .io_config(SBMux_C72_N24254_O_3_C_5_io_config),
    .io_out(SBMux_C72_N24254_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C72_N24254_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C72_N24254_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C72_N24254_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C72_N24254_O_3_C_5_io_arst)
  );
  MuxNInput_O0_C4_SCAOptSB SBMux_C76_N24256_O_0_C_4 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C76_N24256_O_0_C_4_io_in),
    .io_config(SBMux_C76_N24256_O_0_C_4_io_config),
    .io_out(SBMux_C76_N24256_O_0_C_4_io_out),
    .io_loopBreak(SBMux_C76_N24256_O_0_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C76_N24256_O_0_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C76_N24256_O_0_C_4_io_cnstClk),
    .io_arst(SBMux_C76_N24256_O_0_C_4_io_arst)
  );
  MuxNInput_O4_C6_SCAOptSB SBMux_C1_N28731_O_4_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C1_N28731_O_4_C_6_io_in),
    .io_config(SBMux_C1_N28731_O_4_C_6_io_config),
    .io_out(SBMux_C1_N28731_O_4_C_6_io_out),
    .io_loopBreak(SBMux_C1_N28731_O_4_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C1_N28731_O_4_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C1_N28731_O_4_C_6_io_cnstClk),
    .io_arst(SBMux_C1_N28731_O_4_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C9_N28739_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C9_N28739_O_3_C_6_io_in),
    .io_config(SBMux_C9_N28739_O_3_C_6_io_config),
    .io_out(SBMux_C9_N28739_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C9_N28739_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C9_N28739_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C9_N28739_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C9_N28739_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C17_N28747_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C17_N28747_O_3_C_5_io_in),
    .io_config(SBMux_C17_N28747_O_3_C_5_io_config),
    .io_out(SBMux_C17_N28747_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C17_N28747_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C17_N28747_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C17_N28747_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C17_N28747_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C25_N28755_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C25_N28755_O_3_C_5_io_in),
    .io_config(SBMux_C25_N28755_O_3_C_5_io_config),
    .io_out(SBMux_C25_N28755_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C25_N28755_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C25_N28755_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C25_N28755_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C25_N28755_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C33_N28763_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C33_N28763_O_3_C_5_io_in),
    .io_config(SBMux_C33_N28763_O_3_C_5_io_config),
    .io_out(SBMux_C33_N28763_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C33_N28763_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C33_N28763_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C33_N28763_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C33_N28763_O_3_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C41_N28771_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C41_N28771_O_4_C_5_io_in),
    .io_config(SBMux_C41_N28771_O_4_C_5_io_config),
    .io_out(SBMux_C41_N28771_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C41_N28771_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C41_N28771_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C41_N28771_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C41_N28771_O_4_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C49_N28779_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C49_N28779_O_3_C_5_io_in),
    .io_config(SBMux_C49_N28779_O_3_C_5_io_config),
    .io_out(SBMux_C49_N28779_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C49_N28779_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C49_N28779_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C49_N28779_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C49_N28779_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C57_N28787_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C57_N28787_O_3_C_5_io_in),
    .io_config(SBMux_C57_N28787_O_3_C_5_io_config),
    .io_out(SBMux_C57_N28787_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C57_N28787_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C57_N28787_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C57_N28787_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C57_N28787_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C65_N28795_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C65_N28795_O_3_C_5_io_in),
    .io_config(SBMux_C65_N28795_O_3_C_5_io_config),
    .io_out(SBMux_C65_N28795_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C65_N28795_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C65_N28795_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C65_N28795_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C65_N28795_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C73_N28803_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C73_N28803_O_3_C_5_io_in),
    .io_config(SBMux_C73_N28803_O_3_C_5_io_config),
    .io_out(SBMux_C73_N28803_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C73_N28803_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C73_N28803_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C73_N28803_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C73_N28803_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C77_N28829_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C77_N28829_O_3_C_5_io_in),
    .io_config(SBMux_C77_N28829_O_3_C_5_io_config),
    .io_out(SBMux_C77_N28829_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C77_N28829_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C77_N28829_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C77_N28829_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C77_N28829_O_3_C_5_io_arst)
  );
  MuxNInput_O4_C7_SCAOptSB SBMux_C0_N28850_O_4_C_7 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C0_N28850_O_4_C_7_io_in),
    .io_config(SBMux_C0_N28850_O_4_C_7_io_config),
    .io_out(SBMux_C0_N28850_O_4_C_7_io_out),
    .io_loopBreak(SBMux_C0_N28850_O_4_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C0_N28850_O_4_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C0_N28850_O_4_C_7_io_cnstClk),
    .io_arst(SBMux_C0_N28850_O_4_C_7_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C8_N28852_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C8_N28852_O_3_C_6_io_in),
    .io_config(SBMux_C8_N28852_O_3_C_6_io_config),
    .io_out(SBMux_C8_N28852_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C8_N28852_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C8_N28852_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C8_N28852_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C8_N28852_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C16_N28854_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C16_N28854_O_3_C_5_io_in),
    .io_config(SBMux_C16_N28854_O_3_C_5_io_config),
    .io_out(SBMux_C16_N28854_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C16_N28854_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C16_N28854_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C16_N28854_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C16_N28854_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C24_N28856_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C24_N28856_O_3_C_5_io_in),
    .io_config(SBMux_C24_N28856_O_3_C_5_io_config),
    .io_out(SBMux_C24_N28856_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C24_N28856_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C24_N28856_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C24_N28856_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C24_N28856_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C32_N28858_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C32_N28858_O_3_C_5_io_in),
    .io_config(SBMux_C32_N28858_O_3_C_5_io_config),
    .io_out(SBMux_C32_N28858_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C32_N28858_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C32_N28858_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C32_N28858_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C32_N28858_O_3_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C40_N28860_O_4_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C40_N28860_O_4_C_5_io_in),
    .io_config(SBMux_C40_N28860_O_4_C_5_io_config),
    .io_out(SBMux_C40_N28860_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C40_N28860_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C40_N28860_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C40_N28860_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C40_N28860_O_4_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C48_N28862_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C48_N28862_O_3_C_5_io_in),
    .io_config(SBMux_C48_N28862_O_3_C_5_io_config),
    .io_out(SBMux_C48_N28862_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C48_N28862_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C48_N28862_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C48_N28862_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C48_N28862_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C56_N28864_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C56_N28864_O_3_C_5_io_in),
    .io_config(SBMux_C56_N28864_O_3_C_5_io_config),
    .io_out(SBMux_C56_N28864_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C56_N28864_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C56_N28864_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C56_N28864_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C56_N28864_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C64_N28866_O_3_C_5 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C64_N28866_O_3_C_5_io_in),
    .io_config(SBMux_C64_N28866_O_3_C_5_io_config),
    .io_out(SBMux_C64_N28866_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C64_N28866_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C64_N28866_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C64_N28866_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C64_N28866_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C72_N28868_O_3_C_6 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C72_N28868_O_3_C_6_io_in),
    .io_config(SBMux_C72_N28868_O_3_C_6_io_config),
    .io_out(SBMux_C72_N28868_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C72_N28868_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C72_N28868_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C72_N28868_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C72_N28868_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C7_SCAOptSB SBMux_C76_N28870_O_3_C_7 ( // @[TileFull.scala 134:27]
    .io_in(SBMux_C76_N28870_O_3_C_7_io_in),
    .io_config(SBMux_C76_N28870_O_3_C_7_io_config),
    .io_out(SBMux_C76_N28870_O_3_C_7_io_out),
    .io_loopBreak(SBMux_C76_N28870_O_3_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C76_N28870_O_3_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C76_N28870_O_3_C_7_io_cnstClk),
    .io_arst(SBMux_C76_N28870_O_3_C_7_io_arst)
  );
  assign OUT_CHANX_N24242_24 = SBMux_C24_N24242_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24250_56 = SBMux_C56_N24250_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24159_25 = SBMux_C25_N24159_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28868_72 = SBMux_C72_N28868_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28771_41 = SBMux_C41_N28771_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28747_17 = SBMux_C17_N28747_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28858_32 = SBMux_C32_N28858_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19855_45 = logicBlock_OPIN_45; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N28866_64 = SBMux_C64_N28866_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28829_77 = SBMux_C77_N28829_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19861_51 = logicBlock_OPIN_51; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24171_73 = SBMux_C73_N24171_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24155_9 = SBMux_C9_N24155_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24161_33 = SBMux_C33_N24161_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24246_40 = SBMux_C40_N24246_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24165_49 = SBMux_C49_N24165_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24153_1 = SBMux_C1_N24153_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19860_50 = logicBlock_OPIN_50; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24244_32 = SBMux_C32_N24244_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19858_48 = logicBlock_OPIN_48; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24163_41 = SBMux_C41_N24163_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28739_9 = SBMux_C9_N28739_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19864_54 = logicBlock_OPIN_54; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N28860_40 = SBMux_C40_N28860_O_4_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28864_56 = SBMux_C56_N28864_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28850_0 = SBMux_C0_N28850_O_4_C_7_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28755_25 = SBMux_C25_N28755_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28731_1 = SBMux_C1_N28731_O_4_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19865_55 = logicBlock_OPIN_55; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24252_64 = SBMux_C64_N24252_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28870_76 = SBMux_C76_N28870_O_3_C_7_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28795_65 = SBMux_C65_N28795_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28856_24 = SBMux_C24_N28856_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24240_16 = SBMux_C16_N24240_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24238_8 = SBMux_C8_N24238_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19854_44 = logicBlock_OPIN_44; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N28862_48 = SBMux_C48_N28862_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19851_41 = logicBlock_OPIN_41; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24215_77 = SBMux_C77_N24215_O_0_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24256_76 = SBMux_C76_N24256_O_0_C_4_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19853_43 = logicBlock_OPIN_43; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24254_72 = SBMux_C72_N24254_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24248_48 = SBMux_C48_N24248_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19857_47 = logicBlock_OPIN_47; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N28779_49 = SBMux_C49_N28779_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19856_46 = logicBlock_OPIN_46; // @[TileFull.scala 196:12]
  assign OUT_CHANX_N24236_0 = SBMux_C0_N24236_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19863_53 = logicBlock_OPIN_53; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N28854_16 = SBMux_C16_N28854_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19859_49 = logicBlock_OPIN_49; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N28803_73 = SBMux_C73_N28803_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24167_57 = SBMux_C57_N24167_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19866_56 = logicBlock_OPIN_56; // @[TileFull.scala 196:12]
  assign OUT_OPIN_N19852_42 = logicBlock_OPIN_42; // @[TileFull.scala 196:12]
  assign OUT_CHANY_N28763_33 = SBMux_C33_N28763_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24157_17 = SBMux_C17_N24157_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28852_8 = SBMux_C8_N28852_O_3_C_6_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANX_N24169_65 = SBMux_C65_N24169_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_CHANY_N28787_57 = SBMux_C57_N28787_O_3_C_5_io_out; // @[TileFull.scala 138:23]
  assign OUT_OPIN_N19862_52 = logicBlock_OPIN_52; // @[TileFull.scala 196:12]
  assign ioConf_confOut = configBlock_ioBundle_confOut; // @[TileFull.scala 73:12]
  assign ioConf_scan_out = configBlock_ioBundle_scan_out; // @[TileFull.scala 73:12]
  assign logicBlock_IPIN_0 = CBMux_IPIN0_N19810_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_1 = CBMux_IPIN1_N19811_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_2 = CBMux_IPIN2_N19812_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_3 = CBMux_IPIN3_N19813_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_4 = CBMux_IPIN4_N19814_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_5 = CBMux_IPIN5_N19815_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_6 = CBMux_IPIN6_N19816_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_7 = CBMux_IPIN7_N19817_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_8 = CBMux_IPIN8_N19818_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_9 = CBMux_IPIN9_N19819_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_10 = CBMux_IPIN10_N19820_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_11 = CBMux_IPIN11_N19821_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_12 = CBMux_IPIN12_N19822_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_13 = CBMux_IPIN13_N19823_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_14 = CBMux_IPIN14_N19824_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_15 = CBMux_IPIN15_N19825_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_16 = CBMux_IPIN16_N19826_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_17 = CBMux_IPIN17_N19827_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_18 = CBMux_IPIN18_N19828_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_19 = CBMux_IPIN19_N19829_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_20 = CBMux_IPIN20_N19830_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_21 = CBMux_IPIN21_N19831_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_22 = CBMux_IPIN22_N19832_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_23 = CBMux_IPIN23_N19833_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_24 = CBMux_IPIN24_N19834_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_25 = CBMux_IPIN25_N19835_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_26 = CBMux_IPIN26_N19836_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_27 = CBMux_IPIN27_N19837_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_28 = CBMux_IPIN28_N19838_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_29 = CBMux_IPIN29_N19839_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_30 = CBMux_IPIN30_N19840_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_IPIN_31 = CBMux_IPIN31_N19841_io_out; // @[TileFull.scala 100:42]
  assign logicBlock_clock = clock; // @[TileFull.scala 192:26]
  assign logicBlock_reset = reset; // @[TileFull.scala 193:26]
  assign logicBlock_ioPad_i = ioPad_i[15:0]; // @[TileFull.scala 202:32]
  assign logicBlock_configBits = configBlock_ioBundle_confOut[161:0]; // @[TileFull.scala 191:31]
  assign logicBlock_gndLBouts = ctrlSignals_gndBlkOuts; // @[TileFull.scala 189:30]
  assign configBlock_clock = ctrlSignals_confClock; // @[TileFull.scala 74:27]
  assign configBlock_ioBundle_scan_in = ioConf_scan_in; // @[TileFull.scala 73:12]
  assign configBlock_ioBundle_scan_en = ioConf_scan_en; // @[TileFull.scala 73:12]
  assign CBMux_IPIN0_N19810_io_in = {CBMux_IPIN0_N19810_io_in_hi,CBMux_IPIN0_N19810_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN0_N19810_io_config = configBlock_ioBundle_confOut[164:161]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN0_N19810_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN0_N19810_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN0_N19810_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN1_N19811_io_in = {CBMux_IPIN1_N19811_io_in_hi,CBMux_IPIN1_N19811_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN1_N19811_io_config = configBlock_ioBundle_confOut[168:165]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN1_N19811_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN1_N19811_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN1_N19811_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN2_N19812_io_in = {CBMux_IPIN2_N19812_io_in_hi,CBMux_IPIN2_N19812_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN2_N19812_io_config = configBlock_ioBundle_confOut[172:169]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN2_N19812_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN2_N19812_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN2_N19812_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN3_N19813_io_in = {CBMux_IPIN3_N19813_io_in_hi,CBMux_IPIN3_N19813_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN3_N19813_io_config = configBlock_ioBundle_confOut[176:173]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN3_N19813_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN3_N19813_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN3_N19813_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN4_N19814_io_in = {CBMux_IPIN4_N19814_io_in_hi,CBMux_IPIN4_N19814_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN4_N19814_io_config = configBlock_ioBundle_confOut[180:177]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN4_N19814_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN4_N19814_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN4_N19814_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN5_N19815_io_in = {CBMux_IPIN5_N19815_io_in_hi,CBMux_IPIN5_N19815_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN5_N19815_io_config = configBlock_ioBundle_confOut[184:181]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN5_N19815_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN5_N19815_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN5_N19815_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN6_N19816_io_in = {CBMux_IPIN6_N19816_io_in_hi,CBMux_IPIN6_N19816_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN6_N19816_io_config = configBlock_ioBundle_confOut[188:185]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN6_N19816_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN6_N19816_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN6_N19816_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN7_N19817_io_in = {CBMux_IPIN7_N19817_io_in_hi,CBMux_IPIN7_N19817_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN7_N19817_io_config = configBlock_ioBundle_confOut[192:189]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN7_N19817_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN7_N19817_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN7_N19817_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN8_N19818_io_in = {CBMux_IPIN8_N19818_io_in_hi,CBMux_IPIN8_N19818_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN8_N19818_io_config = configBlock_ioBundle_confOut[196:193]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN8_N19818_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN8_N19818_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN8_N19818_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN9_N19819_io_in = {CBMux_IPIN9_N19819_io_in_hi,CBMux_IPIN9_N19819_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN9_N19819_io_config = configBlock_ioBundle_confOut[200:197]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN9_N19819_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN9_N19819_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN9_N19819_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN10_N19820_io_in = {CBMux_IPIN10_N19820_io_in_hi,CBMux_IPIN10_N19820_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN10_N19820_io_config = configBlock_ioBundle_confOut[204:201]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN10_N19820_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN10_N19820_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN10_N19820_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN11_N19821_io_in = {CBMux_IPIN11_N19821_io_in_hi,CBMux_IPIN11_N19821_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN11_N19821_io_config = configBlock_ioBundle_confOut[208:205]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN11_N19821_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN11_N19821_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN11_N19821_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN12_N19822_io_in = {CBMux_IPIN12_N19822_io_in_hi,CBMux_IPIN12_N19822_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN12_N19822_io_config = configBlock_ioBundle_confOut[212:209]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN12_N19822_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN12_N19822_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN12_N19822_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN13_N19823_io_in = {CBMux_IPIN13_N19823_io_in_hi,CBMux_IPIN13_N19823_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN13_N19823_io_config = configBlock_ioBundle_confOut[216:213]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN13_N19823_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN13_N19823_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN13_N19823_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN14_N19824_io_in = {CBMux_IPIN14_N19824_io_in_hi,CBMux_IPIN14_N19824_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN14_N19824_io_config = configBlock_ioBundle_confOut[220:217]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN14_N19824_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN14_N19824_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN14_N19824_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN15_N19825_io_in = {CBMux_IPIN15_N19825_io_in_hi,CBMux_IPIN15_N19825_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN15_N19825_io_config = configBlock_ioBundle_confOut[224:221]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN15_N19825_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN15_N19825_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN15_N19825_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN16_N19826_io_in = {CBMux_IPIN16_N19826_io_in_hi,CBMux_IPIN16_N19826_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN16_N19826_io_config = configBlock_ioBundle_confOut[228:225]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN16_N19826_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN16_N19826_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN16_N19826_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN17_N19827_io_in = {CBMux_IPIN17_N19827_io_in_hi,CBMux_IPIN17_N19827_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN17_N19827_io_config = configBlock_ioBundle_confOut[232:229]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN17_N19827_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN17_N19827_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN17_N19827_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN18_N19828_io_in = {CBMux_IPIN18_N19828_io_in_hi,CBMux_IPIN18_N19828_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN18_N19828_io_config = configBlock_ioBundle_confOut[236:233]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN18_N19828_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN18_N19828_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN18_N19828_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN19_N19829_io_in = {CBMux_IPIN19_N19829_io_in_hi,CBMux_IPIN19_N19829_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN19_N19829_io_config = configBlock_ioBundle_confOut[240:237]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN19_N19829_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN19_N19829_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN19_N19829_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN20_N19830_io_in = {CBMux_IPIN20_N19830_io_in_hi,CBMux_IPIN20_N19830_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN20_N19830_io_config = configBlock_ioBundle_confOut[244:241]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN20_N19830_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN20_N19830_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN20_N19830_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN21_N19831_io_in = {CBMux_IPIN21_N19831_io_in_hi,CBMux_IPIN21_N19831_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN21_N19831_io_config = configBlock_ioBundle_confOut[248:245]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN21_N19831_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN21_N19831_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN21_N19831_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN22_N19832_io_in = {CBMux_IPIN22_N19832_io_in_hi,CBMux_IPIN22_N19832_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN22_N19832_io_config = configBlock_ioBundle_confOut[252:249]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN22_N19832_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN22_N19832_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN22_N19832_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN23_N19833_io_in = {CBMux_IPIN23_N19833_io_in_hi,CBMux_IPIN23_N19833_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN23_N19833_io_config = configBlock_ioBundle_confOut[256:253]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN23_N19833_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN23_N19833_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN23_N19833_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN24_N19834_io_in = {CBMux_IPIN24_N19834_io_in_hi,CBMux_IPIN24_N19834_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN24_N19834_io_config = configBlock_ioBundle_confOut[260:257]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN24_N19834_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN24_N19834_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN24_N19834_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN25_N19835_io_in = {CBMux_IPIN25_N19835_io_in_hi,CBMux_IPIN25_N19835_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN25_N19835_io_config = configBlock_ioBundle_confOut[264:261]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN25_N19835_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN25_N19835_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN25_N19835_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN26_N19836_io_in = {CBMux_IPIN26_N19836_io_in_hi,CBMux_IPIN26_N19836_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN26_N19836_io_config = configBlock_ioBundle_confOut[268:265]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN26_N19836_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN26_N19836_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN26_N19836_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN27_N19837_io_in = {CBMux_IPIN27_N19837_io_in_hi,CBMux_IPIN27_N19837_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN27_N19837_io_config = configBlock_ioBundle_confOut[272:269]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN27_N19837_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN27_N19837_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN27_N19837_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN28_N19838_io_in = {CBMux_IPIN28_N19838_io_in_hi,CBMux_IPIN22_N19832_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN28_N19838_io_config = configBlock_ioBundle_confOut[276:273]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN28_N19838_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN28_N19838_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN28_N19838_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN29_N19839_io_in = {CBMux_IPIN29_N19839_io_in_hi,CBMux_IPIN29_N19839_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN29_N19839_io_config = configBlock_ioBundle_confOut[280:277]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN29_N19839_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN29_N19839_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN29_N19839_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN30_N19840_io_in = {CBMux_IPIN30_N19840_io_in_hi,CBMux_IPIN18_N19828_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN30_N19840_io_config = configBlock_ioBundle_confOut[284:281]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN30_N19840_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN30_N19840_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN30_N19840_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN31_N19841_io_in = {CBMux_IPIN31_N19841_io_in_hi,CBMux_IPIN31_N19841_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN31_N19841_io_config = configBlock_ioBundle_confOut[288:285]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN31_N19841_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN31_N19841_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN31_N19841_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN32_N19842_io_in = {CBMux_IPIN32_N19842_io_in_hi,CBMux_IPIN32_N19842_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN32_N19842_io_config = configBlock_ioBundle_confOut[292:289]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN32_N19842_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN32_N19842_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN32_N19842_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN33_N19843_io_in = {CBMux_IPIN33_N19843_io_in_hi,CBMux_IPIN33_N19843_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN33_N19843_io_config = configBlock_ioBundle_confOut[296:293]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN33_N19843_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN33_N19843_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN33_N19843_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN34_N19844_io_in = {CBMux_IPIN34_N19844_io_in_hi,CBMux_IPIN34_N19844_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN34_N19844_io_config = configBlock_ioBundle_confOut[300:297]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN34_N19844_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN34_N19844_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN34_N19844_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN35_N19845_io_in = {CBMux_IPIN34_N19844_io_in_hi,CBMux_IPIN34_N19844_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN35_N19845_io_config = configBlock_ioBundle_confOut[304:301]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN35_N19845_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN35_N19845_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN35_N19845_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN36_N19846_io_in = {CBMux_IPIN36_N19846_io_in_hi,CBMux_IPIN36_N19846_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN36_N19846_io_config = configBlock_ioBundle_confOut[308:305]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN36_N19846_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN36_N19846_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN36_N19846_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN37_N19847_io_in = {CBMux_IPIN37_N19847_io_in_hi,CBMux_IPIN37_N19847_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN37_N19847_io_config = configBlock_ioBundle_confOut[312:309]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN37_N19847_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN37_N19847_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN37_N19847_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN38_N19848_io_in = {CBMux_IPIN38_N19848_io_in_hi,CBMux_IPIN38_N19848_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN38_N19848_io_config = configBlock_ioBundle_confOut[316:313]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN38_N19848_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN38_N19848_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN38_N19848_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign CBMux_IPIN39_N19849_io_in = {CBMux_IPIN33_N19843_io_in_hi,CBMux_IPIN33_N19843_io_in_lo}; // @[TileFull.scala 166:8]
  assign CBMux_IPIN39_N19849_io_config = configBlock_ioBundle_confOut[320:317]; // @[TileFull.scala 104:60]
  assign CBMux_IPIN39_N19849_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 107:28]
  assign CBMux_IPIN39_N19849_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 108:26]
  assign CBMux_IPIN39_N19849_io_arst = ctrlSignals_arst; // @[TileFull.scala 109:23]
  assign SBMux_C1_N24153_O_3_C_6_io_in = {SBMux_C1_N24153_O_3_C_6_io_in_hi,SBMux_C1_N24153_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C1_N24153_O_3_C_6_io_config = configBlock_ioBundle_confOut[324:321]; // @[TileFull.scala 142:60]
  assign SBMux_C1_N24153_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C1_N24153_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C1_N24153_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C1_N24153_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C9_N24155_O_3_C_6_io_in = {SBMux_C9_N24155_O_3_C_6_io_in_hi,SBMux_C9_N24155_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C9_N24155_O_3_C_6_io_config = configBlock_ioBundle_confOut[328:325]; // @[TileFull.scala 142:60]
  assign SBMux_C9_N24155_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C9_N24155_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C9_N24155_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C9_N24155_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C17_N24157_O_3_C_6_io_in = {SBMux_C17_N24157_O_3_C_6_io_in_hi,SBMux_C17_N24157_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C17_N24157_O_3_C_6_io_config = configBlock_ioBundle_confOut[332:329]; // @[TileFull.scala 142:60]
  assign SBMux_C17_N24157_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C17_N24157_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C17_N24157_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C17_N24157_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C25_N24159_O_3_C_6_io_in = {SBMux_C25_N24159_O_3_C_6_io_in_hi,SBMux_C25_N24159_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C25_N24159_O_3_C_6_io_config = configBlock_ioBundle_confOut[336:333]; // @[TileFull.scala 142:60]
  assign SBMux_C25_N24159_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C25_N24159_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C25_N24159_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C25_N24159_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C33_N24161_O_3_C_5_io_in = {SBMux_C33_N24161_O_3_C_5_io_in_hi,SBMux_C33_N24161_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C33_N24161_O_3_C_5_io_config = configBlock_ioBundle_confOut[340:337]; // @[TileFull.scala 142:60]
  assign SBMux_C33_N24161_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C33_N24161_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C33_N24161_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C33_N24161_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C41_N24163_O_3_C_5_io_in = {SBMux_C41_N24163_O_3_C_5_io_in_hi,SBMux_C41_N24163_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C41_N24163_O_3_C_5_io_config = configBlock_ioBundle_confOut[344:341]; // @[TileFull.scala 142:60]
  assign SBMux_C41_N24163_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C41_N24163_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C41_N24163_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C41_N24163_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C49_N24165_O_3_C_5_io_in = {SBMux_C49_N24165_O_3_C_5_io_in_hi,SBMux_C49_N24165_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C49_N24165_O_3_C_5_io_config = configBlock_ioBundle_confOut[348:345]; // @[TileFull.scala 142:60]
  assign SBMux_C49_N24165_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C49_N24165_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C49_N24165_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C49_N24165_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C57_N24167_O_3_C_5_io_in = {SBMux_C57_N24167_O_3_C_5_io_in_hi,SBMux_C57_N24167_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C57_N24167_O_3_C_5_io_config = configBlock_ioBundle_confOut[352:349]; // @[TileFull.scala 142:60]
  assign SBMux_C57_N24167_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C57_N24167_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C57_N24167_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C57_N24167_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C65_N24169_O_3_C_5_io_in = {SBMux_C65_N24169_O_3_C_5_io_in_hi,SBMux_C65_N24169_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C65_N24169_O_3_C_5_io_config = configBlock_ioBundle_confOut[356:353]; // @[TileFull.scala 142:60]
  assign SBMux_C65_N24169_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C65_N24169_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C65_N24169_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C65_N24169_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C73_N24171_O_3_C_6_io_in = {SBMux_C73_N24171_O_3_C_6_io_in_hi,SBMux_C73_N24171_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C73_N24171_O_3_C_6_io_config = configBlock_ioBundle_confOut[360:357]; // @[TileFull.scala 142:60]
  assign SBMux_C73_N24171_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C73_N24171_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C73_N24171_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C73_N24171_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C77_N24215_O_0_C_6_io_in = {SBMux_C77_N24215_O_0_C_6_io_in_hi,SBMux_C77_N24215_O_0_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C77_N24215_O_0_C_6_io_config = configBlock_ioBundle_confOut[364:361]; // @[TileFull.scala 142:60]
  assign SBMux_C77_N24215_O_0_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C77_N24215_O_0_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C77_N24215_O_0_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C77_N24215_O_0_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C0_N24236_O_3_C_5_io_in = {SBMux_C0_N24236_O_3_C_5_io_in_hi,SBMux_C0_N24236_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C0_N24236_O_3_C_5_io_config = configBlock_ioBundle_confOut[368:365]; // @[TileFull.scala 142:60]
  assign SBMux_C0_N24236_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C0_N24236_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C0_N24236_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C0_N24236_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C8_N24238_O_3_C_6_io_in = {SBMux_C8_N24238_O_3_C_6_io_in_hi,SBMux_C8_N24238_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C8_N24238_O_3_C_6_io_config = configBlock_ioBundle_confOut[372:369]; // @[TileFull.scala 142:60]
  assign SBMux_C8_N24238_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C8_N24238_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C8_N24238_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C8_N24238_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C16_N24240_O_3_C_6_io_in = {SBMux_C16_N24240_O_3_C_6_io_in_hi,SBMux_C16_N24240_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C16_N24240_O_3_C_6_io_config = configBlock_ioBundle_confOut[376:373]; // @[TileFull.scala 142:60]
  assign SBMux_C16_N24240_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C16_N24240_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C16_N24240_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C16_N24240_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C24_N24242_O_3_C_6_io_in = {SBMux_C24_N24242_O_3_C_6_io_in_hi,SBMux_C24_N24242_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C24_N24242_O_3_C_6_io_config = configBlock_ioBundle_confOut[380:377]; // @[TileFull.scala 142:60]
  assign SBMux_C24_N24242_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C24_N24242_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C24_N24242_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C24_N24242_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C32_N24244_O_3_C_5_io_in = {SBMux_C32_N24244_O_3_C_5_io_in_hi,SBMux_C32_N24244_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C32_N24244_O_3_C_5_io_config = configBlock_ioBundle_confOut[384:381]; // @[TileFull.scala 142:60]
  assign SBMux_C32_N24244_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C32_N24244_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C32_N24244_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C32_N24244_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C40_N24246_O_3_C_5_io_in = {SBMux_C40_N24246_O_3_C_5_io_in_hi,SBMux_C40_N24246_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C40_N24246_O_3_C_5_io_config = configBlock_ioBundle_confOut[388:385]; // @[TileFull.scala 142:60]
  assign SBMux_C40_N24246_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C40_N24246_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C40_N24246_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C40_N24246_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C48_N24248_O_3_C_5_io_in = {SBMux_C48_N24248_O_3_C_5_io_in_hi,SBMux_C48_N24248_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C48_N24248_O_3_C_5_io_config = configBlock_ioBundle_confOut[392:389]; // @[TileFull.scala 142:60]
  assign SBMux_C48_N24248_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C48_N24248_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C48_N24248_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C48_N24248_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C56_N24250_O_3_C_5_io_in = {SBMux_C56_N24250_O_3_C_5_io_in_hi,SBMux_C56_N24250_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C56_N24250_O_3_C_5_io_config = configBlock_ioBundle_confOut[396:393]; // @[TileFull.scala 142:60]
  assign SBMux_C56_N24250_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C56_N24250_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C56_N24250_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C56_N24250_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C64_N24252_O_3_C_5_io_in = {SBMux_C64_N24252_O_3_C_5_io_in_hi,SBMux_C64_N24252_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C64_N24252_O_3_C_5_io_config = configBlock_ioBundle_confOut[400:397]; // @[TileFull.scala 142:60]
  assign SBMux_C64_N24252_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C64_N24252_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C64_N24252_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C64_N24252_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C72_N24254_O_3_C_5_io_in = {SBMux_C72_N24254_O_3_C_5_io_in_hi,SBMux_C72_N24254_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C72_N24254_O_3_C_5_io_config = configBlock_ioBundle_confOut[404:401]; // @[TileFull.scala 142:60]
  assign SBMux_C72_N24254_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C72_N24254_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C72_N24254_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C72_N24254_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C76_N24256_O_0_C_4_io_in = {SBMux_C76_N24256_O_0_C_4_io_in_hi,SBMux_C76_N24256_O_0_C_4_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C76_N24256_O_0_C_4_io_config = configBlock_ioBundle_confOut[407:405]; // @[TileFull.scala 142:60]
  assign SBMux_C76_N24256_O_0_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C76_N24256_O_0_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C76_N24256_O_0_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C76_N24256_O_0_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C1_N28731_O_4_C_6_io_in = {SBMux_C1_N28731_O_4_C_6_io_in_hi,SBMux_C1_N28731_O_4_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C1_N28731_O_4_C_6_io_config = configBlock_ioBundle_confOut[411:408]; // @[TileFull.scala 142:60]
  assign SBMux_C1_N28731_O_4_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C1_N28731_O_4_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C1_N28731_O_4_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C1_N28731_O_4_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C9_N28739_O_3_C_6_io_in = {SBMux_C9_N28739_O_3_C_6_io_in_hi,SBMux_C9_N28739_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C9_N28739_O_3_C_6_io_config = configBlock_ioBundle_confOut[415:412]; // @[TileFull.scala 142:60]
  assign SBMux_C9_N28739_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C9_N28739_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C9_N28739_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C9_N28739_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C17_N28747_O_3_C_5_io_in = {SBMux_C17_N28747_O_3_C_5_io_in_hi,SBMux_C17_N28747_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C17_N28747_O_3_C_5_io_config = configBlock_ioBundle_confOut[419:416]; // @[TileFull.scala 142:60]
  assign SBMux_C17_N28747_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C17_N28747_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C17_N28747_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C17_N28747_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C25_N28755_O_3_C_5_io_in = {SBMux_C25_N28755_O_3_C_5_io_in_hi,SBMux_C25_N28755_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C25_N28755_O_3_C_5_io_config = configBlock_ioBundle_confOut[423:420]; // @[TileFull.scala 142:60]
  assign SBMux_C25_N28755_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C25_N28755_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C25_N28755_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C25_N28755_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C33_N28763_O_3_C_5_io_in = {SBMux_C33_N28763_O_3_C_5_io_in_hi,SBMux_C33_N28763_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C33_N28763_O_3_C_5_io_config = configBlock_ioBundle_confOut[427:424]; // @[TileFull.scala 142:60]
  assign SBMux_C33_N28763_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C33_N28763_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C33_N28763_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C33_N28763_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C41_N28771_O_4_C_5_io_in = {SBMux_C41_N28771_O_4_C_5_io_in_hi,SBMux_C41_N28771_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C41_N28771_O_4_C_5_io_config = configBlock_ioBundle_confOut[431:428]; // @[TileFull.scala 142:60]
  assign SBMux_C41_N28771_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C41_N28771_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C41_N28771_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C41_N28771_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C49_N28779_O_3_C_5_io_in = {SBMux_C49_N28779_O_3_C_5_io_in_hi,SBMux_C49_N28779_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C49_N28779_O_3_C_5_io_config = configBlock_ioBundle_confOut[435:432]; // @[TileFull.scala 142:60]
  assign SBMux_C49_N28779_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C49_N28779_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C49_N28779_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C49_N28779_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C57_N28787_O_3_C_5_io_in = {SBMux_C57_N28787_O_3_C_5_io_in_hi,SBMux_C57_N28787_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C57_N28787_O_3_C_5_io_config = configBlock_ioBundle_confOut[439:436]; // @[TileFull.scala 142:60]
  assign SBMux_C57_N28787_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C57_N28787_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C57_N28787_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C57_N28787_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C65_N28795_O_3_C_5_io_in = {SBMux_C65_N28795_O_3_C_5_io_in_hi,SBMux_C65_N28795_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C65_N28795_O_3_C_5_io_config = configBlock_ioBundle_confOut[443:440]; // @[TileFull.scala 142:60]
  assign SBMux_C65_N28795_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C65_N28795_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C65_N28795_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C65_N28795_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C73_N28803_O_3_C_5_io_in = {SBMux_C73_N28803_O_3_C_5_io_in_hi,SBMux_C73_N28803_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C73_N28803_O_3_C_5_io_config = configBlock_ioBundle_confOut[447:444]; // @[TileFull.scala 142:60]
  assign SBMux_C73_N28803_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C73_N28803_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C73_N28803_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C73_N28803_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C77_N28829_O_3_C_5_io_in = {SBMux_C77_N28829_O_3_C_5_io_in_hi,SBMux_C77_N28829_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C77_N28829_O_3_C_5_io_config = configBlock_ioBundle_confOut[451:448]; // @[TileFull.scala 142:60]
  assign SBMux_C77_N28829_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C77_N28829_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C77_N28829_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C77_N28829_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C0_N28850_O_4_C_7_io_in = {SBMux_C0_N28850_O_4_C_7_io_in_hi,SBMux_C0_N28850_O_4_C_7_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C0_N28850_O_4_C_7_io_config = configBlock_ioBundle_confOut[455:452]; // @[TileFull.scala 142:60]
  assign SBMux_C0_N28850_O_4_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C0_N28850_O_4_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C0_N28850_O_4_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C0_N28850_O_4_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C8_N28852_O_3_C_6_io_in = {SBMux_C8_N28852_O_3_C_6_io_in_hi,SBMux_C8_N28852_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C8_N28852_O_3_C_6_io_config = configBlock_ioBundle_confOut[459:456]; // @[TileFull.scala 142:60]
  assign SBMux_C8_N28852_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C8_N28852_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C8_N28852_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C8_N28852_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C16_N28854_O_3_C_5_io_in = {SBMux_C16_N28854_O_3_C_5_io_in_hi,SBMux_C16_N28854_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C16_N28854_O_3_C_5_io_config = configBlock_ioBundle_confOut[463:460]; // @[TileFull.scala 142:60]
  assign SBMux_C16_N28854_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C16_N28854_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C16_N28854_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C16_N28854_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C24_N28856_O_3_C_5_io_in = {SBMux_C24_N28856_O_3_C_5_io_in_hi,SBMux_C24_N28856_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C24_N28856_O_3_C_5_io_config = configBlock_ioBundle_confOut[467:464]; // @[TileFull.scala 142:60]
  assign SBMux_C24_N28856_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C24_N28856_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C24_N28856_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C24_N28856_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C32_N28858_O_3_C_5_io_in = {SBMux_C32_N28858_O_3_C_5_io_in_hi,SBMux_C32_N28858_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C32_N28858_O_3_C_5_io_config = configBlock_ioBundle_confOut[471:468]; // @[TileFull.scala 142:60]
  assign SBMux_C32_N28858_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C32_N28858_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C32_N28858_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C32_N28858_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C40_N28860_O_4_C_5_io_in = {SBMux_C40_N28860_O_4_C_5_io_in_hi,SBMux_C40_N28860_O_4_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C40_N28860_O_4_C_5_io_config = configBlock_ioBundle_confOut[475:472]; // @[TileFull.scala 142:60]
  assign SBMux_C40_N28860_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C40_N28860_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C40_N28860_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C40_N28860_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C48_N28862_O_3_C_5_io_in = {SBMux_C48_N28862_O_3_C_5_io_in_hi,SBMux_C48_N28862_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C48_N28862_O_3_C_5_io_config = configBlock_ioBundle_confOut[479:476]; // @[TileFull.scala 142:60]
  assign SBMux_C48_N28862_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C48_N28862_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C48_N28862_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C48_N28862_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C56_N28864_O_3_C_5_io_in = {SBMux_C56_N28864_O_3_C_5_io_in_hi,SBMux_C56_N28864_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C56_N28864_O_3_C_5_io_config = configBlock_ioBundle_confOut[483:480]; // @[TileFull.scala 142:60]
  assign SBMux_C56_N28864_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C56_N28864_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C56_N28864_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C56_N28864_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C64_N28866_O_3_C_5_io_in = {SBMux_C64_N28866_O_3_C_5_io_in_hi,SBMux_C64_N28866_O_3_C_5_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C64_N28866_O_3_C_5_io_config = configBlock_ioBundle_confOut[487:484]; // @[TileFull.scala 142:60]
  assign SBMux_C64_N28866_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C64_N28866_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C64_N28866_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C64_N28866_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C72_N28868_O_3_C_6_io_in = {SBMux_C72_N28868_O_3_C_6_io_in_hi,SBMux_C72_N28868_O_3_C_6_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C72_N28868_O_3_C_6_io_config = configBlock_ioBundle_confOut[491:488]; // @[TileFull.scala 142:60]
  assign SBMux_C72_N28868_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C72_N28868_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C72_N28868_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C72_N28868_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
  assign SBMux_C76_N28870_O_3_C_7_io_in = {SBMux_C76_N28870_O_3_C_7_io_in_hi,SBMux_C76_N28870_O_3_C_7_io_in_lo}; // @[TileFull.scala 183:11]
  assign SBMux_C76_N28870_O_3_C_7_io_config = configBlock_ioBundle_confOut[495:492]; // @[TileFull.scala 142:60]
  assign SBMux_C76_N28870_O_3_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 146:28]
  assign SBMux_C76_N28870_O_3_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 149:27]
  assign SBMux_C76_N28870_O_3_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 147:26]
  assign SBMux_C76_N28870_O_3_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 148:23]
endmodule
