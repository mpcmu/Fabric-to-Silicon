//module  \$_DFF_PN0_ (input D, C, R, output Q); ARL0DFF _TECHMAP_REPLACE_ (.D(D), .Q(Q), .C(C), .R(R)); wire _TECHMAP_REMOVEINIT_Q_ = 1; endmodule
//module  \$_DFF_PN1_ (input D, C, R, output Q); ARL1DFF _TECHMAP_REPLACE_ (.D(D), .Q(Q), .C(C), .R(R)); wire _TECHMAP_REMOVEINIT_Q_ = 1; endmodule
//module  \$_DFF_P (input D, C, R, output Q); R0DFF _TECHMAP_REPLACE_ (.D(D), .Q(Q), .C(C), .R(R)); wire _TECHMAP_REMOVEINIT_Q_ = 1; endmodule
//module  \$_DFF_PN1_ (input D, C, R, output Q); ARL1DFF _TECHMAP_REPLACE_ (.D(D), .Q(Q), .C(C), .R(R)); wire _TECHMAP_REMOVEINIT_Q_ = 1; endmodule
