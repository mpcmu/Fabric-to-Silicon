module BUFx2_ASAP7_75t_L (A, Y);
	input A;
	output Y;
	assign Y = A;
endmodule
