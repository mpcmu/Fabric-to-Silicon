module ScanConf_Tile_7_3_clbalutile(
  input          clock,
  input          reset,
  output [511:0] ioBundle_confOut,
  input  [15:0]  ioBundle_scan_in,
  input          ioBundle_scan_en,
  output [15:0]  ioBundle_scan_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
`endif // RANDOMIZE_REG_INIT
  reg  confReg_0; // @[ScanConf.scala 32:20]
  reg  confReg_1; // @[ScanConf.scala 32:20]
  reg  confReg_2; // @[ScanConf.scala 32:20]
  reg  confReg_3; // @[ScanConf.scala 32:20]
  reg  confReg_4; // @[ScanConf.scala 32:20]
  reg  confReg_5; // @[ScanConf.scala 32:20]
  reg  confReg_6; // @[ScanConf.scala 32:20]
  reg  confReg_7; // @[ScanConf.scala 32:20]
  reg  confReg_8; // @[ScanConf.scala 32:20]
  reg  confReg_9; // @[ScanConf.scala 32:20]
  reg  confReg_10; // @[ScanConf.scala 32:20]
  reg  confReg_11; // @[ScanConf.scala 32:20]
  reg  confReg_12; // @[ScanConf.scala 32:20]
  reg  confReg_13; // @[ScanConf.scala 32:20]
  reg  confReg_14; // @[ScanConf.scala 32:20]
  reg  confReg_15; // @[ScanConf.scala 32:20]
  reg  confReg_16; // @[ScanConf.scala 32:20]
  reg  confReg_17; // @[ScanConf.scala 32:20]
  reg  confReg_18; // @[ScanConf.scala 32:20]
  reg  confReg_19; // @[ScanConf.scala 32:20]
  reg  confReg_20; // @[ScanConf.scala 32:20]
  reg  confReg_21; // @[ScanConf.scala 32:20]
  reg  confReg_22; // @[ScanConf.scala 32:20]
  reg  confReg_23; // @[ScanConf.scala 32:20]
  reg  confReg_24; // @[ScanConf.scala 32:20]
  reg  confReg_25; // @[ScanConf.scala 32:20]
  reg  confReg_26; // @[ScanConf.scala 32:20]
  reg  confReg_27; // @[ScanConf.scala 32:20]
  reg  confReg_28; // @[ScanConf.scala 32:20]
  reg  confReg_29; // @[ScanConf.scala 32:20]
  reg  confReg_30; // @[ScanConf.scala 32:20]
  reg  confReg_31; // @[ScanConf.scala 32:20]
  reg  confReg_32; // @[ScanConf.scala 32:20]
  reg  confReg_33; // @[ScanConf.scala 32:20]
  reg  confReg_34; // @[ScanConf.scala 32:20]
  reg  confReg_35; // @[ScanConf.scala 32:20]
  reg  confReg_36; // @[ScanConf.scala 32:20]
  reg  confReg_37; // @[ScanConf.scala 32:20]
  reg  confReg_38; // @[ScanConf.scala 32:20]
  reg  confReg_39; // @[ScanConf.scala 32:20]
  reg  confReg_40; // @[ScanConf.scala 32:20]
  reg  confReg_41; // @[ScanConf.scala 32:20]
  reg  confReg_42; // @[ScanConf.scala 32:20]
  reg  confReg_43; // @[ScanConf.scala 32:20]
  reg  confReg_44; // @[ScanConf.scala 32:20]
  reg  confReg_45; // @[ScanConf.scala 32:20]
  reg  confReg_46; // @[ScanConf.scala 32:20]
  reg  confReg_47; // @[ScanConf.scala 32:20]
  reg  confReg_48; // @[ScanConf.scala 32:20]
  reg  confReg_49; // @[ScanConf.scala 32:20]
  reg  confReg_50; // @[ScanConf.scala 32:20]
  reg  confReg_51; // @[ScanConf.scala 32:20]
  reg  confReg_52; // @[ScanConf.scala 32:20]
  reg  confReg_53; // @[ScanConf.scala 32:20]
  reg  confReg_54; // @[ScanConf.scala 32:20]
  reg  confReg_55; // @[ScanConf.scala 32:20]
  reg  confReg_56; // @[ScanConf.scala 32:20]
  reg  confReg_57; // @[ScanConf.scala 32:20]
  reg  confReg_58; // @[ScanConf.scala 32:20]
  reg  confReg_59; // @[ScanConf.scala 32:20]
  reg  confReg_60; // @[ScanConf.scala 32:20]
  reg  confReg_61; // @[ScanConf.scala 32:20]
  reg  confReg_62; // @[ScanConf.scala 32:20]
  reg  confReg_63; // @[ScanConf.scala 32:20]
  reg  confReg_64; // @[ScanConf.scala 32:20]
  reg  confReg_65; // @[ScanConf.scala 32:20]
  reg  confReg_66; // @[ScanConf.scala 32:20]
  reg  confReg_67; // @[ScanConf.scala 32:20]
  reg  confReg_68; // @[ScanConf.scala 32:20]
  reg  confReg_69; // @[ScanConf.scala 32:20]
  reg  confReg_70; // @[ScanConf.scala 32:20]
  reg  confReg_71; // @[ScanConf.scala 32:20]
  reg  confReg_72; // @[ScanConf.scala 32:20]
  reg  confReg_73; // @[ScanConf.scala 32:20]
  reg  confReg_74; // @[ScanConf.scala 32:20]
  reg  confReg_75; // @[ScanConf.scala 32:20]
  reg  confReg_76; // @[ScanConf.scala 32:20]
  reg  confReg_77; // @[ScanConf.scala 32:20]
  reg  confReg_78; // @[ScanConf.scala 32:20]
  reg  confReg_79; // @[ScanConf.scala 32:20]
  reg  confReg_80; // @[ScanConf.scala 32:20]
  reg  confReg_81; // @[ScanConf.scala 32:20]
  reg  confReg_82; // @[ScanConf.scala 32:20]
  reg  confReg_83; // @[ScanConf.scala 32:20]
  reg  confReg_84; // @[ScanConf.scala 32:20]
  reg  confReg_85; // @[ScanConf.scala 32:20]
  reg  confReg_86; // @[ScanConf.scala 32:20]
  reg  confReg_87; // @[ScanConf.scala 32:20]
  reg  confReg_88; // @[ScanConf.scala 32:20]
  reg  confReg_89; // @[ScanConf.scala 32:20]
  reg  confReg_90; // @[ScanConf.scala 32:20]
  reg  confReg_91; // @[ScanConf.scala 32:20]
  reg  confReg_92; // @[ScanConf.scala 32:20]
  reg  confReg_93; // @[ScanConf.scala 32:20]
  reg  confReg_94; // @[ScanConf.scala 32:20]
  reg  confReg_95; // @[ScanConf.scala 32:20]
  reg  confReg_96; // @[ScanConf.scala 32:20]
  reg  confReg_97; // @[ScanConf.scala 32:20]
  reg  confReg_98; // @[ScanConf.scala 32:20]
  reg  confReg_99; // @[ScanConf.scala 32:20]
  reg  confReg_100; // @[ScanConf.scala 32:20]
  reg  confReg_101; // @[ScanConf.scala 32:20]
  reg  confReg_102; // @[ScanConf.scala 32:20]
  reg  confReg_103; // @[ScanConf.scala 32:20]
  reg  confReg_104; // @[ScanConf.scala 32:20]
  reg  confReg_105; // @[ScanConf.scala 32:20]
  reg  confReg_106; // @[ScanConf.scala 32:20]
  reg  confReg_107; // @[ScanConf.scala 32:20]
  reg  confReg_108; // @[ScanConf.scala 32:20]
  reg  confReg_109; // @[ScanConf.scala 32:20]
  reg  confReg_110; // @[ScanConf.scala 32:20]
  reg  confReg_111; // @[ScanConf.scala 32:20]
  reg  confReg_112; // @[ScanConf.scala 32:20]
  reg  confReg_113; // @[ScanConf.scala 32:20]
  reg  confReg_114; // @[ScanConf.scala 32:20]
  reg  confReg_115; // @[ScanConf.scala 32:20]
  reg  confReg_116; // @[ScanConf.scala 32:20]
  reg  confReg_117; // @[ScanConf.scala 32:20]
  reg  confReg_118; // @[ScanConf.scala 32:20]
  reg  confReg_119; // @[ScanConf.scala 32:20]
  reg  confReg_120; // @[ScanConf.scala 32:20]
  reg  confReg_121; // @[ScanConf.scala 32:20]
  reg  confReg_122; // @[ScanConf.scala 32:20]
  reg  confReg_123; // @[ScanConf.scala 32:20]
  reg  confReg_124; // @[ScanConf.scala 32:20]
  reg  confReg_125; // @[ScanConf.scala 32:20]
  reg  confReg_126; // @[ScanConf.scala 32:20]
  reg  confReg_127; // @[ScanConf.scala 32:20]
  reg  confReg_128; // @[ScanConf.scala 32:20]
  reg  confReg_129; // @[ScanConf.scala 32:20]
  reg  confReg_130; // @[ScanConf.scala 32:20]
  reg  confReg_131; // @[ScanConf.scala 32:20]
  reg  confReg_132; // @[ScanConf.scala 32:20]
  reg  confReg_133; // @[ScanConf.scala 32:20]
  reg  confReg_134; // @[ScanConf.scala 32:20]
  reg  confReg_135; // @[ScanConf.scala 32:20]
  reg  confReg_136; // @[ScanConf.scala 32:20]
  reg  confReg_137; // @[ScanConf.scala 32:20]
  reg  confReg_138; // @[ScanConf.scala 32:20]
  reg  confReg_139; // @[ScanConf.scala 32:20]
  reg  confReg_140; // @[ScanConf.scala 32:20]
  reg  confReg_141; // @[ScanConf.scala 32:20]
  reg  confReg_142; // @[ScanConf.scala 32:20]
  reg  confReg_143; // @[ScanConf.scala 32:20]
  reg  confReg_144; // @[ScanConf.scala 32:20]
  reg  confReg_145; // @[ScanConf.scala 32:20]
  reg  confReg_146; // @[ScanConf.scala 32:20]
  reg  confReg_147; // @[ScanConf.scala 32:20]
  reg  confReg_148; // @[ScanConf.scala 32:20]
  reg  confReg_149; // @[ScanConf.scala 32:20]
  reg  confReg_150; // @[ScanConf.scala 32:20]
  reg  confReg_151; // @[ScanConf.scala 32:20]
  reg  confReg_152; // @[ScanConf.scala 32:20]
  reg  confReg_153; // @[ScanConf.scala 32:20]
  reg  confReg_154; // @[ScanConf.scala 32:20]
  reg  confReg_155; // @[ScanConf.scala 32:20]
  reg  confReg_156; // @[ScanConf.scala 32:20]
  reg  confReg_157; // @[ScanConf.scala 32:20]
  reg  confReg_158; // @[ScanConf.scala 32:20]
  reg  confReg_159; // @[ScanConf.scala 32:20]
  reg  confReg_160; // @[ScanConf.scala 32:20]
  reg  confReg_161; // @[ScanConf.scala 32:20]
  reg  confReg_162; // @[ScanConf.scala 32:20]
  reg  confReg_163; // @[ScanConf.scala 32:20]
  reg  confReg_164; // @[ScanConf.scala 32:20]
  reg  confReg_165; // @[ScanConf.scala 32:20]
  reg  confReg_166; // @[ScanConf.scala 32:20]
  reg  confReg_167; // @[ScanConf.scala 32:20]
  reg  confReg_168; // @[ScanConf.scala 32:20]
  reg  confReg_169; // @[ScanConf.scala 32:20]
  reg  confReg_170; // @[ScanConf.scala 32:20]
  reg  confReg_171; // @[ScanConf.scala 32:20]
  reg  confReg_172; // @[ScanConf.scala 32:20]
  reg  confReg_173; // @[ScanConf.scala 32:20]
  reg  confReg_174; // @[ScanConf.scala 32:20]
  reg  confReg_175; // @[ScanConf.scala 32:20]
  reg  confReg_176; // @[ScanConf.scala 32:20]
  reg  confReg_177; // @[ScanConf.scala 32:20]
  reg  confReg_178; // @[ScanConf.scala 32:20]
  reg  confReg_179; // @[ScanConf.scala 32:20]
  reg  confReg_180; // @[ScanConf.scala 32:20]
  reg  confReg_181; // @[ScanConf.scala 32:20]
  reg  confReg_182; // @[ScanConf.scala 32:20]
  reg  confReg_183; // @[ScanConf.scala 32:20]
  reg  confReg_184; // @[ScanConf.scala 32:20]
  reg  confReg_185; // @[ScanConf.scala 32:20]
  reg  confReg_186; // @[ScanConf.scala 32:20]
  reg  confReg_187; // @[ScanConf.scala 32:20]
  reg  confReg_188; // @[ScanConf.scala 32:20]
  reg  confReg_189; // @[ScanConf.scala 32:20]
  reg  confReg_190; // @[ScanConf.scala 32:20]
  reg  confReg_191; // @[ScanConf.scala 32:20]
  reg  confReg_192; // @[ScanConf.scala 32:20]
  reg  confReg_193; // @[ScanConf.scala 32:20]
  reg  confReg_194; // @[ScanConf.scala 32:20]
  reg  confReg_195; // @[ScanConf.scala 32:20]
  reg  confReg_196; // @[ScanConf.scala 32:20]
  reg  confReg_197; // @[ScanConf.scala 32:20]
  reg  confReg_198; // @[ScanConf.scala 32:20]
  reg  confReg_199; // @[ScanConf.scala 32:20]
  reg  confReg_200; // @[ScanConf.scala 32:20]
  reg  confReg_201; // @[ScanConf.scala 32:20]
  reg  confReg_202; // @[ScanConf.scala 32:20]
  reg  confReg_203; // @[ScanConf.scala 32:20]
  reg  confReg_204; // @[ScanConf.scala 32:20]
  reg  confReg_205; // @[ScanConf.scala 32:20]
  reg  confReg_206; // @[ScanConf.scala 32:20]
  reg  confReg_207; // @[ScanConf.scala 32:20]
  reg  confReg_208; // @[ScanConf.scala 32:20]
  reg  confReg_209; // @[ScanConf.scala 32:20]
  reg  confReg_210; // @[ScanConf.scala 32:20]
  reg  confReg_211; // @[ScanConf.scala 32:20]
  reg  confReg_212; // @[ScanConf.scala 32:20]
  reg  confReg_213; // @[ScanConf.scala 32:20]
  reg  confReg_214; // @[ScanConf.scala 32:20]
  reg  confReg_215; // @[ScanConf.scala 32:20]
  reg  confReg_216; // @[ScanConf.scala 32:20]
  reg  confReg_217; // @[ScanConf.scala 32:20]
  reg  confReg_218; // @[ScanConf.scala 32:20]
  reg  confReg_219; // @[ScanConf.scala 32:20]
  reg  confReg_220; // @[ScanConf.scala 32:20]
  reg  confReg_221; // @[ScanConf.scala 32:20]
  reg  confReg_222; // @[ScanConf.scala 32:20]
  reg  confReg_223; // @[ScanConf.scala 32:20]
  reg  confReg_224; // @[ScanConf.scala 32:20]
  reg  confReg_225; // @[ScanConf.scala 32:20]
  reg  confReg_226; // @[ScanConf.scala 32:20]
  reg  confReg_227; // @[ScanConf.scala 32:20]
  reg  confReg_228; // @[ScanConf.scala 32:20]
  reg  confReg_229; // @[ScanConf.scala 32:20]
  reg  confReg_230; // @[ScanConf.scala 32:20]
  reg  confReg_231; // @[ScanConf.scala 32:20]
  reg  confReg_232; // @[ScanConf.scala 32:20]
  reg  confReg_233; // @[ScanConf.scala 32:20]
  reg  confReg_234; // @[ScanConf.scala 32:20]
  reg  confReg_235; // @[ScanConf.scala 32:20]
  reg  confReg_236; // @[ScanConf.scala 32:20]
  reg  confReg_237; // @[ScanConf.scala 32:20]
  reg  confReg_238; // @[ScanConf.scala 32:20]
  reg  confReg_239; // @[ScanConf.scala 32:20]
  reg  confReg_240; // @[ScanConf.scala 32:20]
  reg  confReg_241; // @[ScanConf.scala 32:20]
  reg  confReg_242; // @[ScanConf.scala 32:20]
  reg  confReg_243; // @[ScanConf.scala 32:20]
  reg  confReg_244; // @[ScanConf.scala 32:20]
  reg  confReg_245; // @[ScanConf.scala 32:20]
  reg  confReg_246; // @[ScanConf.scala 32:20]
  reg  confReg_247; // @[ScanConf.scala 32:20]
  reg  confReg_248; // @[ScanConf.scala 32:20]
  reg  confReg_249; // @[ScanConf.scala 32:20]
  reg  confReg_250; // @[ScanConf.scala 32:20]
  reg  confReg_251; // @[ScanConf.scala 32:20]
  reg  confReg_252; // @[ScanConf.scala 32:20]
  reg  confReg_253; // @[ScanConf.scala 32:20]
  reg  confReg_254; // @[ScanConf.scala 32:20]
  reg  confReg_255; // @[ScanConf.scala 32:20]
  reg  confReg_256; // @[ScanConf.scala 32:20]
  reg  confReg_257; // @[ScanConf.scala 32:20]
  reg  confReg_258; // @[ScanConf.scala 32:20]
  reg  confReg_259; // @[ScanConf.scala 32:20]
  reg  confReg_260; // @[ScanConf.scala 32:20]
  reg  confReg_261; // @[ScanConf.scala 32:20]
  reg  confReg_262; // @[ScanConf.scala 32:20]
  reg  confReg_263; // @[ScanConf.scala 32:20]
  reg  confReg_264; // @[ScanConf.scala 32:20]
  reg  confReg_265; // @[ScanConf.scala 32:20]
  reg  confReg_266; // @[ScanConf.scala 32:20]
  reg  confReg_267; // @[ScanConf.scala 32:20]
  reg  confReg_268; // @[ScanConf.scala 32:20]
  reg  confReg_269; // @[ScanConf.scala 32:20]
  reg  confReg_270; // @[ScanConf.scala 32:20]
  reg  confReg_271; // @[ScanConf.scala 32:20]
  reg  confReg_272; // @[ScanConf.scala 32:20]
  reg  confReg_273; // @[ScanConf.scala 32:20]
  reg  confReg_274; // @[ScanConf.scala 32:20]
  reg  confReg_275; // @[ScanConf.scala 32:20]
  reg  confReg_276; // @[ScanConf.scala 32:20]
  reg  confReg_277; // @[ScanConf.scala 32:20]
  reg  confReg_278; // @[ScanConf.scala 32:20]
  reg  confReg_279; // @[ScanConf.scala 32:20]
  reg  confReg_280; // @[ScanConf.scala 32:20]
  reg  confReg_281; // @[ScanConf.scala 32:20]
  reg  confReg_282; // @[ScanConf.scala 32:20]
  reg  confReg_283; // @[ScanConf.scala 32:20]
  reg  confReg_284; // @[ScanConf.scala 32:20]
  reg  confReg_285; // @[ScanConf.scala 32:20]
  reg  confReg_286; // @[ScanConf.scala 32:20]
  reg  confReg_287; // @[ScanConf.scala 32:20]
  reg  confReg_288; // @[ScanConf.scala 32:20]
  reg  confReg_289; // @[ScanConf.scala 32:20]
  reg  confReg_290; // @[ScanConf.scala 32:20]
  reg  confReg_291; // @[ScanConf.scala 32:20]
  reg  confReg_292; // @[ScanConf.scala 32:20]
  reg  confReg_293; // @[ScanConf.scala 32:20]
  reg  confReg_294; // @[ScanConf.scala 32:20]
  reg  confReg_295; // @[ScanConf.scala 32:20]
  reg  confReg_296; // @[ScanConf.scala 32:20]
  reg  confReg_297; // @[ScanConf.scala 32:20]
  reg  confReg_298; // @[ScanConf.scala 32:20]
  reg  confReg_299; // @[ScanConf.scala 32:20]
  reg  confReg_300; // @[ScanConf.scala 32:20]
  reg  confReg_301; // @[ScanConf.scala 32:20]
  reg  confReg_302; // @[ScanConf.scala 32:20]
  reg  confReg_303; // @[ScanConf.scala 32:20]
  reg  confReg_304; // @[ScanConf.scala 32:20]
  reg  confReg_305; // @[ScanConf.scala 32:20]
  reg  confReg_306; // @[ScanConf.scala 32:20]
  reg  confReg_307; // @[ScanConf.scala 32:20]
  reg  confReg_308; // @[ScanConf.scala 32:20]
  reg  confReg_309; // @[ScanConf.scala 32:20]
  reg  confReg_310; // @[ScanConf.scala 32:20]
  reg  confReg_311; // @[ScanConf.scala 32:20]
  reg  confReg_312; // @[ScanConf.scala 32:20]
  reg  confReg_313; // @[ScanConf.scala 32:20]
  reg  confReg_314; // @[ScanConf.scala 32:20]
  reg  confReg_315; // @[ScanConf.scala 32:20]
  reg  confReg_316; // @[ScanConf.scala 32:20]
  reg  confReg_317; // @[ScanConf.scala 32:20]
  reg  confReg_318; // @[ScanConf.scala 32:20]
  reg  confReg_319; // @[ScanConf.scala 32:20]
  reg  confReg_320; // @[ScanConf.scala 32:20]
  reg  confReg_321; // @[ScanConf.scala 32:20]
  reg  confReg_322; // @[ScanConf.scala 32:20]
  reg  confReg_323; // @[ScanConf.scala 32:20]
  reg  confReg_324; // @[ScanConf.scala 32:20]
  reg  confReg_325; // @[ScanConf.scala 32:20]
  reg  confReg_326; // @[ScanConf.scala 32:20]
  reg  confReg_327; // @[ScanConf.scala 32:20]
  reg  confReg_328; // @[ScanConf.scala 32:20]
  reg  confReg_329; // @[ScanConf.scala 32:20]
  reg  confReg_330; // @[ScanConf.scala 32:20]
  reg  confReg_331; // @[ScanConf.scala 32:20]
  reg  confReg_332; // @[ScanConf.scala 32:20]
  reg  confReg_333; // @[ScanConf.scala 32:20]
  reg  confReg_334; // @[ScanConf.scala 32:20]
  reg  confReg_335; // @[ScanConf.scala 32:20]
  reg  confReg_336; // @[ScanConf.scala 32:20]
  reg  confReg_337; // @[ScanConf.scala 32:20]
  reg  confReg_338; // @[ScanConf.scala 32:20]
  reg  confReg_339; // @[ScanConf.scala 32:20]
  reg  confReg_340; // @[ScanConf.scala 32:20]
  reg  confReg_341; // @[ScanConf.scala 32:20]
  reg  confReg_342; // @[ScanConf.scala 32:20]
  reg  confReg_343; // @[ScanConf.scala 32:20]
  reg  confReg_344; // @[ScanConf.scala 32:20]
  reg  confReg_345; // @[ScanConf.scala 32:20]
  reg  confReg_346; // @[ScanConf.scala 32:20]
  reg  confReg_347; // @[ScanConf.scala 32:20]
  reg  confReg_348; // @[ScanConf.scala 32:20]
  reg  confReg_349; // @[ScanConf.scala 32:20]
  reg  confReg_350; // @[ScanConf.scala 32:20]
  reg  confReg_351; // @[ScanConf.scala 32:20]
  reg  confReg_352; // @[ScanConf.scala 32:20]
  reg  confReg_353; // @[ScanConf.scala 32:20]
  reg  confReg_354; // @[ScanConf.scala 32:20]
  reg  confReg_355; // @[ScanConf.scala 32:20]
  reg  confReg_356; // @[ScanConf.scala 32:20]
  reg  confReg_357; // @[ScanConf.scala 32:20]
  reg  confReg_358; // @[ScanConf.scala 32:20]
  reg  confReg_359; // @[ScanConf.scala 32:20]
  reg  confReg_360; // @[ScanConf.scala 32:20]
  reg  confReg_361; // @[ScanConf.scala 32:20]
  reg  confReg_362; // @[ScanConf.scala 32:20]
  reg  confReg_363; // @[ScanConf.scala 32:20]
  reg  confReg_364; // @[ScanConf.scala 32:20]
  reg  confReg_365; // @[ScanConf.scala 32:20]
  reg  confReg_366; // @[ScanConf.scala 32:20]
  reg  confReg_367; // @[ScanConf.scala 32:20]
  reg  confReg_368; // @[ScanConf.scala 32:20]
  reg  confReg_369; // @[ScanConf.scala 32:20]
  reg  confReg_370; // @[ScanConf.scala 32:20]
  reg  confReg_371; // @[ScanConf.scala 32:20]
  reg  confReg_372; // @[ScanConf.scala 32:20]
  reg  confReg_373; // @[ScanConf.scala 32:20]
  reg  confReg_374; // @[ScanConf.scala 32:20]
  reg  confReg_375; // @[ScanConf.scala 32:20]
  reg  confReg_376; // @[ScanConf.scala 32:20]
  reg  confReg_377; // @[ScanConf.scala 32:20]
  reg  confReg_378; // @[ScanConf.scala 32:20]
  reg  confReg_379; // @[ScanConf.scala 32:20]
  reg  confReg_380; // @[ScanConf.scala 32:20]
  reg  confReg_381; // @[ScanConf.scala 32:20]
  reg  confReg_382; // @[ScanConf.scala 32:20]
  reg  confReg_383; // @[ScanConf.scala 32:20]
  reg  confReg_384; // @[ScanConf.scala 32:20]
  reg  confReg_385; // @[ScanConf.scala 32:20]
  reg  confReg_386; // @[ScanConf.scala 32:20]
  reg  confReg_387; // @[ScanConf.scala 32:20]
  reg  confReg_388; // @[ScanConf.scala 32:20]
  reg  confReg_389; // @[ScanConf.scala 32:20]
  reg  confReg_390; // @[ScanConf.scala 32:20]
  reg  confReg_391; // @[ScanConf.scala 32:20]
  reg  confReg_392; // @[ScanConf.scala 32:20]
  reg  confReg_393; // @[ScanConf.scala 32:20]
  reg  confReg_394; // @[ScanConf.scala 32:20]
  reg  confReg_395; // @[ScanConf.scala 32:20]
  reg  confReg_396; // @[ScanConf.scala 32:20]
  reg  confReg_397; // @[ScanConf.scala 32:20]
  reg  confReg_398; // @[ScanConf.scala 32:20]
  reg  confReg_399; // @[ScanConf.scala 32:20]
  reg  confReg_400; // @[ScanConf.scala 32:20]
  reg  confReg_401; // @[ScanConf.scala 32:20]
  reg  confReg_402; // @[ScanConf.scala 32:20]
  reg  confReg_403; // @[ScanConf.scala 32:20]
  reg  confReg_404; // @[ScanConf.scala 32:20]
  reg  confReg_405; // @[ScanConf.scala 32:20]
  reg  confReg_406; // @[ScanConf.scala 32:20]
  reg  confReg_407; // @[ScanConf.scala 32:20]
  reg  confReg_408; // @[ScanConf.scala 32:20]
  reg  confReg_409; // @[ScanConf.scala 32:20]
  reg  confReg_410; // @[ScanConf.scala 32:20]
  reg  confReg_411; // @[ScanConf.scala 32:20]
  reg  confReg_412; // @[ScanConf.scala 32:20]
  reg  confReg_413; // @[ScanConf.scala 32:20]
  reg  confReg_414; // @[ScanConf.scala 32:20]
  reg  confReg_415; // @[ScanConf.scala 32:20]
  reg  confReg_416; // @[ScanConf.scala 32:20]
  reg  confReg_417; // @[ScanConf.scala 32:20]
  reg  confReg_418; // @[ScanConf.scala 32:20]
  reg  confReg_419; // @[ScanConf.scala 32:20]
  reg  confReg_420; // @[ScanConf.scala 32:20]
  reg  confReg_421; // @[ScanConf.scala 32:20]
  reg  confReg_422; // @[ScanConf.scala 32:20]
  reg  confReg_423; // @[ScanConf.scala 32:20]
  reg  confReg_424; // @[ScanConf.scala 32:20]
  reg  confReg_425; // @[ScanConf.scala 32:20]
  reg  confReg_426; // @[ScanConf.scala 32:20]
  reg  confReg_427; // @[ScanConf.scala 32:20]
  reg  confReg_428; // @[ScanConf.scala 32:20]
  reg  confReg_429; // @[ScanConf.scala 32:20]
  reg  confReg_430; // @[ScanConf.scala 32:20]
  reg  confReg_431; // @[ScanConf.scala 32:20]
  reg  confReg_432; // @[ScanConf.scala 32:20]
  reg  confReg_433; // @[ScanConf.scala 32:20]
  reg  confReg_434; // @[ScanConf.scala 32:20]
  reg  confReg_435; // @[ScanConf.scala 32:20]
  reg  confReg_436; // @[ScanConf.scala 32:20]
  reg  confReg_437; // @[ScanConf.scala 32:20]
  reg  confReg_438; // @[ScanConf.scala 32:20]
  reg  confReg_439; // @[ScanConf.scala 32:20]
  reg  confReg_440; // @[ScanConf.scala 32:20]
  reg  confReg_441; // @[ScanConf.scala 32:20]
  reg  confReg_442; // @[ScanConf.scala 32:20]
  reg  confReg_443; // @[ScanConf.scala 32:20]
  reg  confReg_444; // @[ScanConf.scala 32:20]
  reg  confReg_445; // @[ScanConf.scala 32:20]
  reg  confReg_446; // @[ScanConf.scala 32:20]
  reg  confReg_447; // @[ScanConf.scala 32:20]
  reg  confReg_448; // @[ScanConf.scala 32:20]
  reg  confReg_449; // @[ScanConf.scala 32:20]
  reg  confReg_450; // @[ScanConf.scala 32:20]
  reg  confReg_451; // @[ScanConf.scala 32:20]
  reg  confReg_452; // @[ScanConf.scala 32:20]
  reg  confReg_453; // @[ScanConf.scala 32:20]
  reg  confReg_454; // @[ScanConf.scala 32:20]
  reg  confReg_455; // @[ScanConf.scala 32:20]
  reg  confReg_456; // @[ScanConf.scala 32:20]
  reg  confReg_457; // @[ScanConf.scala 32:20]
  reg  confReg_458; // @[ScanConf.scala 32:20]
  reg  confReg_459; // @[ScanConf.scala 32:20]
  reg  confReg_460; // @[ScanConf.scala 32:20]
  reg  confReg_461; // @[ScanConf.scala 32:20]
  reg  confReg_462; // @[ScanConf.scala 32:20]
  reg  confReg_463; // @[ScanConf.scala 32:20]
  reg  confReg_464; // @[ScanConf.scala 32:20]
  reg  confReg_465; // @[ScanConf.scala 32:20]
  reg  confReg_466; // @[ScanConf.scala 32:20]
  reg  confReg_467; // @[ScanConf.scala 32:20]
  reg  confReg_468; // @[ScanConf.scala 32:20]
  reg  confReg_469; // @[ScanConf.scala 32:20]
  reg  confReg_470; // @[ScanConf.scala 32:20]
  reg  confReg_471; // @[ScanConf.scala 32:20]
  reg  confReg_472; // @[ScanConf.scala 32:20]
  reg  confReg_473; // @[ScanConf.scala 32:20]
  reg  confReg_474; // @[ScanConf.scala 32:20]
  reg  confReg_475; // @[ScanConf.scala 32:20]
  reg  confReg_476; // @[ScanConf.scala 32:20]
  reg  confReg_477; // @[ScanConf.scala 32:20]
  reg  confReg_478; // @[ScanConf.scala 32:20]
  reg  confReg_479; // @[ScanConf.scala 32:20]
  reg  confReg_480; // @[ScanConf.scala 32:20]
  reg  confReg_481; // @[ScanConf.scala 32:20]
  reg  confReg_482; // @[ScanConf.scala 32:20]
  reg  confReg_483; // @[ScanConf.scala 32:20]
  reg  confReg_484; // @[ScanConf.scala 32:20]
  reg  confReg_485; // @[ScanConf.scala 32:20]
  reg  confReg_486; // @[ScanConf.scala 32:20]
  reg  confReg_487; // @[ScanConf.scala 32:20]
  reg  confReg_488; // @[ScanConf.scala 32:20]
  reg  confReg_489; // @[ScanConf.scala 32:20]
  reg  confReg_490; // @[ScanConf.scala 32:20]
  reg  confReg_491; // @[ScanConf.scala 32:20]
  reg  confReg_492; // @[ScanConf.scala 32:20]
  reg  confReg_493; // @[ScanConf.scala 32:20]
  reg  confReg_494; // @[ScanConf.scala 32:20]
  reg  confReg_495; // @[ScanConf.scala 32:20]
  reg  confReg_496; // @[ScanConf.scala 32:20]
  reg  confReg_497; // @[ScanConf.scala 32:20]
  reg  confReg_498; // @[ScanConf.scala 32:20]
  reg  confReg_499; // @[ScanConf.scala 32:20]
  reg  confReg_500; // @[ScanConf.scala 32:20]
  reg  confReg_501; // @[ScanConf.scala 32:20]
  reg  confReg_502; // @[ScanConf.scala 32:20]
  reg  confReg_503; // @[ScanConf.scala 32:20]
  reg  confReg_504; // @[ScanConf.scala 32:20]
  reg  confReg_505; // @[ScanConf.scala 32:20]
  reg  confReg_506; // @[ScanConf.scala 32:20]
  reg  confReg_507; // @[ScanConf.scala 32:20]
  reg  confReg_508; // @[ScanConf.scala 32:20]
  reg  confReg_509; // @[ScanConf.scala 32:20]
  reg  confReg_510; // @[ScanConf.scala 32:20]
  reg  confReg_511; // @[ScanConf.scala 32:20]
  wire [7:0] io_scan_out_lo = {confReg_7,confReg_6,confReg_5,confReg_4,confReg_3,confReg_2,confReg_1,confReg_0}; // @[ScanConf.scala 46:47]
  wire [7:0] io_scan_out_hi = {confReg_15,confReg_14,confReg_13,confReg_12,confReg_11,confReg_10,confReg_9,confReg_8}; // @[ScanConf.scala 46:47]
  wire [15:0] io_scan_out = {confReg_15,confReg_14,confReg_13,confReg_12,confReg_11,confReg_10,confReg_9,confReg_8,
    io_scan_out_lo}; // @[ScanConf.scala 46:47]
  wire [7:0] io_confOut_lo_lo_lo_lo_hi_lo = {confReg_23,confReg_22,confReg_21,confReg_20,confReg_19,confReg_18,
    confReg_17,confReg_16}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_lo_lo_lo = {confReg_31,confReg_30,confReg_29,confReg_28,confReg_27,confReg_26,confReg_25,
    confReg_24,io_confOut_lo_lo_lo_lo_hi_lo,io_scan_out}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_lo_hi_lo_lo = {confReg_39,confReg_38,confReg_37,confReg_36,confReg_35,confReg_34,
    confReg_33,confReg_32}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_lo_lo_hi_lo = {confReg_47,confReg_46,confReg_45,confReg_44,confReg_43,confReg_42,confReg_41,
    confReg_40,io_confOut_lo_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_lo_hi_hi_lo = {confReg_55,confReg_54,confReg_53,confReg_52,confReg_51,confReg_50,
    confReg_49,confReg_48}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_lo_lo_hi = {confReg_63,confReg_62,confReg_61,confReg_60,confReg_59,confReg_58,confReg_57,
    confReg_56,io_confOut_lo_lo_lo_hi_hi_lo,io_confOut_lo_lo_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_hi_lo_lo_lo = {confReg_71,confReg_70,confReg_69,confReg_68,confReg_67,confReg_66,
    confReg_65,confReg_64}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_lo_hi_lo_lo = {confReg_79,confReg_78,confReg_77,confReg_76,confReg_75,confReg_74,confReg_73,
    confReg_72,io_confOut_lo_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_hi_lo_hi_lo = {confReg_87,confReg_86,confReg_85,confReg_84,confReg_83,confReg_82,
    confReg_81,confReg_80}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_lo_hi_lo = {confReg_95,confReg_94,confReg_93,confReg_92,confReg_91,confReg_90,confReg_89,
    confReg_88,io_confOut_lo_lo_hi_lo_hi_lo,io_confOut_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_hi_hi_lo_lo = {confReg_103,confReg_102,confReg_101,confReg_100,confReg_99,confReg_98,
    confReg_97,confReg_96}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_lo_hi_hi_lo = {confReg_111,confReg_110,confReg_109,confReg_108,confReg_107,confReg_106,
    confReg_105,confReg_104,io_confOut_lo_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_lo_hi_hi_hi_lo = {confReg_119,confReg_118,confReg_117,confReg_116,confReg_115,confReg_114,
    confReg_113,confReg_112}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_lo_hi_hi = {confReg_127,confReg_126,confReg_125,confReg_124,confReg_123,confReg_122,
    confReg_121,confReg_120,io_confOut_lo_lo_hi_hi_hi_lo,io_confOut_lo_lo_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_lo_lo_lo_lo = {confReg_135,confReg_134,confReg_133,confReg_132,confReg_131,confReg_130,
    confReg_129,confReg_128}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_hi_lo_lo_lo = {confReg_143,confReg_142,confReg_141,confReg_140,confReg_139,confReg_138,
    confReg_137,confReg_136,io_confOut_lo_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_lo_lo_hi_lo = {confReg_151,confReg_150,confReg_149,confReg_148,confReg_147,confReg_146,
    confReg_145,confReg_144}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_hi_lo_lo = {confReg_159,confReg_158,confReg_157,confReg_156,confReg_155,confReg_154,
    confReg_153,confReg_152,io_confOut_lo_hi_lo_lo_hi_lo,io_confOut_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_lo_hi_lo_lo = {confReg_167,confReg_166,confReg_165,confReg_164,confReg_163,confReg_162,
    confReg_161,confReg_160}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_hi_lo_hi_lo = {confReg_175,confReg_174,confReg_173,confReg_172,confReg_171,confReg_170,
    confReg_169,confReg_168,io_confOut_lo_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_lo_hi_hi_lo = {confReg_183,confReg_182,confReg_181,confReg_180,confReg_179,confReg_178,
    confReg_177,confReg_176}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_hi_lo_hi = {confReg_191,confReg_190,confReg_189,confReg_188,confReg_187,confReg_186,
    confReg_185,confReg_184,io_confOut_lo_hi_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_hi_lo_lo_lo = {confReg_199,confReg_198,confReg_197,confReg_196,confReg_195,confReg_194,
    confReg_193,confReg_192}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_hi_hi_lo_lo = {confReg_207,confReg_206,confReg_205,confReg_204,confReg_203,confReg_202,
    confReg_201,confReg_200,io_confOut_lo_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_hi_lo_hi_lo = {confReg_215,confReg_214,confReg_213,confReg_212,confReg_211,confReg_210,
    confReg_209,confReg_208}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_hi_hi_lo = {confReg_223,confReg_222,confReg_221,confReg_220,confReg_219,confReg_218,
    confReg_217,confReg_216,io_confOut_lo_hi_hi_lo_hi_lo,io_confOut_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_hi_hi_lo_lo = {confReg_231,confReg_230,confReg_229,confReg_228,confReg_227,confReg_226,
    confReg_225,confReg_224}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_lo_hi_hi_hi_lo = {confReg_239,confReg_238,confReg_237,confReg_236,confReg_235,confReg_234,
    confReg_233,confReg_232,io_confOut_lo_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_lo_hi_hi_hi_hi_lo = {confReg_247,confReg_246,confReg_245,confReg_244,confReg_243,confReg_242,
    confReg_241,confReg_240}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_lo_hi_hi_hi = {confReg_255,confReg_254,confReg_253,confReg_252,confReg_251,confReg_250,
    confReg_249,confReg_248,io_confOut_lo_hi_hi_hi_hi_lo,io_confOut_lo_hi_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [255:0] io_confOut_lo = {io_confOut_lo_hi_hi_hi,io_confOut_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi,
    io_confOut_lo_hi_lo_lo,io_confOut_lo_lo_hi_hi,io_confOut_lo_lo_hi_lo,io_confOut_lo_lo_lo_hi,io_confOut_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_lo_lo_lo_lo = {confReg_263,confReg_262,confReg_261,confReg_260,confReg_259,confReg_258,
    confReg_257,confReg_256}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_lo_lo_lo_lo = {confReg_271,confReg_270,confReg_269,confReg_268,confReg_267,confReg_266,
    confReg_265,confReg_264,io_confOut_hi_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_lo_lo_hi_lo = {confReg_279,confReg_278,confReg_277,confReg_276,confReg_275,confReg_274,
    confReg_273,confReg_272}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_lo_lo_lo = {confReg_287,confReg_286,confReg_285,confReg_284,confReg_283,confReg_282,
    confReg_281,confReg_280,io_confOut_hi_lo_lo_lo_hi_lo,io_confOut_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_lo_hi_lo_lo = {confReg_295,confReg_294,confReg_293,confReg_292,confReg_291,confReg_290,
    confReg_289,confReg_288}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_lo_lo_hi_lo = {confReg_303,confReg_302,confReg_301,confReg_300,confReg_299,confReg_298,
    confReg_297,confReg_296,io_confOut_hi_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_lo_hi_hi_lo = {confReg_311,confReg_310,confReg_309,confReg_308,confReg_307,confReg_306,
    confReg_305,confReg_304}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_lo_lo_hi = {confReg_319,confReg_318,confReg_317,confReg_316,confReg_315,confReg_314,
    confReg_313,confReg_312,io_confOut_hi_lo_lo_hi_hi_lo,io_confOut_hi_lo_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_hi_lo_lo_lo = {confReg_327,confReg_326,confReg_325,confReg_324,confReg_323,confReg_322,
    confReg_321,confReg_320}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_lo_hi_lo_lo = {confReg_335,confReg_334,confReg_333,confReg_332,confReg_331,confReg_330,
    confReg_329,confReg_328,io_confOut_hi_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_hi_lo_hi_lo = {confReg_343,confReg_342,confReg_341,confReg_340,confReg_339,confReg_338,
    confReg_337,confReg_336}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_lo_hi_lo = {confReg_351,confReg_350,confReg_349,confReg_348,confReg_347,confReg_346,
    confReg_345,confReg_344,io_confOut_hi_lo_hi_lo_hi_lo,io_confOut_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_hi_hi_lo_lo = {confReg_359,confReg_358,confReg_357,confReg_356,confReg_355,confReg_354,
    confReg_353,confReg_352}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_lo_hi_hi_lo = {confReg_367,confReg_366,confReg_365,confReg_364,confReg_363,confReg_362,
    confReg_361,confReg_360,io_confOut_hi_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_lo_hi_hi_hi_lo = {confReg_375,confReg_374,confReg_373,confReg_372,confReg_371,confReg_370,
    confReg_369,confReg_368}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_lo_hi_hi = {confReg_383,confReg_382,confReg_381,confReg_380,confReg_379,confReg_378,
    confReg_377,confReg_376,io_confOut_hi_lo_hi_hi_hi_lo,io_confOut_hi_lo_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_lo_lo_lo_lo = {confReg_391,confReg_390,confReg_389,confReg_388,confReg_387,confReg_386,
    confReg_385,confReg_384}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_hi_lo_lo_lo = {confReg_399,confReg_398,confReg_397,confReg_396,confReg_395,confReg_394,
    confReg_393,confReg_392,io_confOut_hi_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_lo_lo_hi_lo = {confReg_407,confReg_406,confReg_405,confReg_404,confReg_403,confReg_402,
    confReg_401,confReg_400}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_hi_lo_lo = {confReg_415,confReg_414,confReg_413,confReg_412,confReg_411,confReg_410,
    confReg_409,confReg_408,io_confOut_hi_hi_lo_lo_hi_lo,io_confOut_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_lo_hi_lo_lo = {confReg_423,confReg_422,confReg_421,confReg_420,confReg_419,confReg_418,
    confReg_417,confReg_416}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_hi_lo_hi_lo = {confReg_431,confReg_430,confReg_429,confReg_428,confReg_427,confReg_426,
    confReg_425,confReg_424,io_confOut_hi_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_lo_hi_hi_lo = {confReg_439,confReg_438,confReg_437,confReg_436,confReg_435,confReg_434,
    confReg_433,confReg_432}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_hi_lo_hi = {confReg_447,confReg_446,confReg_445,confReg_444,confReg_443,confReg_442,
    confReg_441,confReg_440,io_confOut_hi_hi_lo_hi_hi_lo,io_confOut_hi_hi_lo_hi_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_hi_lo_lo_lo = {confReg_455,confReg_454,confReg_453,confReg_452,confReg_451,confReg_450,
    confReg_449,confReg_448}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_hi_hi_lo_lo = {confReg_463,confReg_462,confReg_461,confReg_460,confReg_459,confReg_458,
    confReg_457,confReg_456,io_confOut_hi_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_hi_lo_hi_lo = {confReg_471,confReg_470,confReg_469,confReg_468,confReg_467,confReg_466,
    confReg_465,confReg_464}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_hi_hi_lo = {confReg_479,confReg_478,confReg_477,confReg_476,confReg_475,confReg_474,
    confReg_473,confReg_472,io_confOut_hi_hi_hi_lo_hi_lo,io_confOut_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_hi_hi_lo_lo = {confReg_487,confReg_486,confReg_485,confReg_484,confReg_483,confReg_482,
    confReg_481,confReg_480}; // @[ScanConf.scala 48:25]
  wire [15:0] io_confOut_hi_hi_hi_hi_lo = {confReg_495,confReg_494,confReg_493,confReg_492,confReg_491,confReg_490,
    confReg_489,confReg_488,io_confOut_hi_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [7:0] io_confOut_hi_hi_hi_hi_hi_lo = {confReg_503,confReg_502,confReg_501,confReg_500,confReg_499,confReg_498,
    confReg_497,confReg_496}; // @[ScanConf.scala 48:25]
  wire [31:0] io_confOut_hi_hi_hi_hi = {confReg_511,confReg_510,confReg_509,confReg_508,confReg_507,confReg_506,
    confReg_505,confReg_504,io_confOut_hi_hi_hi_hi_hi_lo,io_confOut_hi_hi_hi_hi_lo}; // @[ScanConf.scala 48:25]
  wire [255:0] io_confOut_hi = {io_confOut_hi_hi_hi_hi,io_confOut_hi_hi_hi_lo,io_confOut_hi_hi_lo_hi,
    io_confOut_hi_hi_lo_lo,io_confOut_hi_lo_hi_hi,io_confOut_hi_lo_hi_lo,io_confOut_hi_lo_lo_hi,io_confOut_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  assign ioBundle_confOut = {io_confOut_hi,io_confOut_lo}; // @[ScanConf.scala 48:25]
  assign ioBundle_scan_out = {io_scan_out_hi,io_scan_out_lo}; // @[ScanConf.scala 46:47]
  always @(posedge clock) begin
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_0 <= confReg_16; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_1 <= confReg_17; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_2 <= confReg_18; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_3 <= confReg_19; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_4 <= confReg_20; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_5 <= confReg_21; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_6 <= confReg_22; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_7 <= confReg_23; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_8 <= confReg_24; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_9 <= confReg_25; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_10 <= confReg_26; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_11 <= confReg_27; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_12 <= confReg_28; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_13 <= confReg_29; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_14 <= confReg_30; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_15 <= confReg_31; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_16 <= confReg_32; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_17 <= confReg_33; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_18 <= confReg_34; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_19 <= confReg_35; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_20 <= confReg_36; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_21 <= confReg_37; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_22 <= confReg_38; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_23 <= confReg_39; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_24 <= confReg_40; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_25 <= confReg_41; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_26 <= confReg_42; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_27 <= confReg_43; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_28 <= confReg_44; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_29 <= confReg_45; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_30 <= confReg_46; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_31 <= confReg_47; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_32 <= confReg_48; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_33 <= confReg_49; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_34 <= confReg_50; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_35 <= confReg_51; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_36 <= confReg_52; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_37 <= confReg_53; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_38 <= confReg_54; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_39 <= confReg_55; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_40 <= confReg_56; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_41 <= confReg_57; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_42 <= confReg_58; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_43 <= confReg_59; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_44 <= confReg_60; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_45 <= confReg_61; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_46 <= confReg_62; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_47 <= confReg_63; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_48 <= confReg_64; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_49 <= confReg_65; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_50 <= confReg_66; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_51 <= confReg_67; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_52 <= confReg_68; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_53 <= confReg_69; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_54 <= confReg_70; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_55 <= confReg_71; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_56 <= confReg_72; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_57 <= confReg_73; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_58 <= confReg_74; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_59 <= confReg_75; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_60 <= confReg_76; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_61 <= confReg_77; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_62 <= confReg_78; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_63 <= confReg_79; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_64 <= confReg_80; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_65 <= confReg_81; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_66 <= confReg_82; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_67 <= confReg_83; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_68 <= confReg_84; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_69 <= confReg_85; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_70 <= confReg_86; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_71 <= confReg_87; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_72 <= confReg_88; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_73 <= confReg_89; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_74 <= confReg_90; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_75 <= confReg_91; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_76 <= confReg_92; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_77 <= confReg_93; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_78 <= confReg_94; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_79 <= confReg_95; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_80 <= confReg_96; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_81 <= confReg_97; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_82 <= confReg_98; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_83 <= confReg_99; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_84 <= confReg_100; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_85 <= confReg_101; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_86 <= confReg_102; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_87 <= confReg_103; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_88 <= confReg_104; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_89 <= confReg_105; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_90 <= confReg_106; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_91 <= confReg_107; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_92 <= confReg_108; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_93 <= confReg_109; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_94 <= confReg_110; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_95 <= confReg_111; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_96 <= confReg_112; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_97 <= confReg_113; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_98 <= confReg_114; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_99 <= confReg_115; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_100 <= confReg_116; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_101 <= confReg_117; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_102 <= confReg_118; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_103 <= confReg_119; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_104 <= confReg_120; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_105 <= confReg_121; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_106 <= confReg_122; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_107 <= confReg_123; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_108 <= confReg_124; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_109 <= confReg_125; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_110 <= confReg_126; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_111 <= confReg_127; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_112 <= confReg_128; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_113 <= confReg_129; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_114 <= confReg_130; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_115 <= confReg_131; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_116 <= confReg_132; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_117 <= confReg_133; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_118 <= confReg_134; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_119 <= confReg_135; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_120 <= confReg_136; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_121 <= confReg_137; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_122 <= confReg_138; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_123 <= confReg_139; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_124 <= confReg_140; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_125 <= confReg_141; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_126 <= confReg_142; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_127 <= confReg_143; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_128 <= confReg_144; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_129 <= confReg_145; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_130 <= confReg_146; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_131 <= confReg_147; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_132 <= confReg_148; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_133 <= confReg_149; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_134 <= confReg_150; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_135 <= confReg_151; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_136 <= confReg_152; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_137 <= confReg_153; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_138 <= confReg_154; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_139 <= confReg_155; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_140 <= confReg_156; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_141 <= confReg_157; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_142 <= confReg_158; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_143 <= confReg_159; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_144 <= confReg_160; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_145 <= confReg_161; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_146 <= confReg_162; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_147 <= confReg_163; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_148 <= confReg_164; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_149 <= confReg_165; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_150 <= confReg_166; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_151 <= confReg_167; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_152 <= confReg_168; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_153 <= confReg_169; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_154 <= confReg_170; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_155 <= confReg_171; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_156 <= confReg_172; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_157 <= confReg_173; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_158 <= confReg_174; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_159 <= confReg_175; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_160 <= confReg_176; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_161 <= confReg_177; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_162 <= confReg_178; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_163 <= confReg_179; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_164 <= confReg_180; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_165 <= confReg_181; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_166 <= confReg_182; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_167 <= confReg_183; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_168 <= confReg_184; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_169 <= confReg_185; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_170 <= confReg_186; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_171 <= confReg_187; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_172 <= confReg_188; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_173 <= confReg_189; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_174 <= confReg_190; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_175 <= confReg_191; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_176 <= confReg_192; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_177 <= confReg_193; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_178 <= confReg_194; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_179 <= confReg_195; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_180 <= confReg_196; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_181 <= confReg_197; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_182 <= confReg_198; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_183 <= confReg_199; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_184 <= confReg_200; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_185 <= confReg_201; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_186 <= confReg_202; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_187 <= confReg_203; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_188 <= confReg_204; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_189 <= confReg_205; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_190 <= confReg_206; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_191 <= confReg_207; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_192 <= confReg_208; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_193 <= confReg_209; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_194 <= confReg_210; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_195 <= confReg_211; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_196 <= confReg_212; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_197 <= confReg_213; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_198 <= confReg_214; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_199 <= confReg_215; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_200 <= confReg_216; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_201 <= confReg_217; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_202 <= confReg_218; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_203 <= confReg_219; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_204 <= confReg_220; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_205 <= confReg_221; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_206 <= confReg_222; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_207 <= confReg_223; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_208 <= confReg_224; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_209 <= confReg_225; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_210 <= confReg_226; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_211 <= confReg_227; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_212 <= confReg_228; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_213 <= confReg_229; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_214 <= confReg_230; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_215 <= confReg_231; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_216 <= confReg_232; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_217 <= confReg_233; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_218 <= confReg_234; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_219 <= confReg_235; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_220 <= confReg_236; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_221 <= confReg_237; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_222 <= confReg_238; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_223 <= confReg_239; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_224 <= confReg_240; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_225 <= confReg_241; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_226 <= confReg_242; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_227 <= confReg_243; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_228 <= confReg_244; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_229 <= confReg_245; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_230 <= confReg_246; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_231 <= confReg_247; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_232 <= confReg_248; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_233 <= confReg_249; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_234 <= confReg_250; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_235 <= confReg_251; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_236 <= confReg_252; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_237 <= confReg_253; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_238 <= confReg_254; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_239 <= confReg_255; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_240 <= confReg_256; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_241 <= confReg_257; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_242 <= confReg_258; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_243 <= confReg_259; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_244 <= confReg_260; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_245 <= confReg_261; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_246 <= confReg_262; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_247 <= confReg_263; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_248 <= confReg_264; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_249 <= confReg_265; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_250 <= confReg_266; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_251 <= confReg_267; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_252 <= confReg_268; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_253 <= confReg_269; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_254 <= confReg_270; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_255 <= confReg_271; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_256 <= confReg_272; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_257 <= confReg_273; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_258 <= confReg_274; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_259 <= confReg_275; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_260 <= confReg_276; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_261 <= confReg_277; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_262 <= confReg_278; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_263 <= confReg_279; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_264 <= confReg_280; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_265 <= confReg_281; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_266 <= confReg_282; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_267 <= confReg_283; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_268 <= confReg_284; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_269 <= confReg_285; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_270 <= confReg_286; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_271 <= confReg_287; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_272 <= confReg_288; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_273 <= confReg_289; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_274 <= confReg_290; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_275 <= confReg_291; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_276 <= confReg_292; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_277 <= confReg_293; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_278 <= confReg_294; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_279 <= confReg_295; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_280 <= confReg_296; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_281 <= confReg_297; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_282 <= confReg_298; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_283 <= confReg_299; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_284 <= confReg_300; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_285 <= confReg_301; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_286 <= confReg_302; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_287 <= confReg_303; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_288 <= confReg_304; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_289 <= confReg_305; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_290 <= confReg_306; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_291 <= confReg_307; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_292 <= confReg_308; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_293 <= confReg_309; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_294 <= confReg_310; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_295 <= confReg_311; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_296 <= confReg_312; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_297 <= confReg_313; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_298 <= confReg_314; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_299 <= confReg_315; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_300 <= confReg_316; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_301 <= confReg_317; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_302 <= confReg_318; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_303 <= confReg_319; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_304 <= confReg_320; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_305 <= confReg_321; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_306 <= confReg_322; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_307 <= confReg_323; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_308 <= confReg_324; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_309 <= confReg_325; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_310 <= confReg_326; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_311 <= confReg_327; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_312 <= confReg_328; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_313 <= confReg_329; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_314 <= confReg_330; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_315 <= confReg_331; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_316 <= confReg_332; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_317 <= confReg_333; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_318 <= confReg_334; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_319 <= confReg_335; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_320 <= confReg_336; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_321 <= confReg_337; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_322 <= confReg_338; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_323 <= confReg_339; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_324 <= confReg_340; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_325 <= confReg_341; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_326 <= confReg_342; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_327 <= confReg_343; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_328 <= confReg_344; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_329 <= confReg_345; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_330 <= confReg_346; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_331 <= confReg_347; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_332 <= confReg_348; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_333 <= confReg_349; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_334 <= confReg_350; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_335 <= confReg_351; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_336 <= confReg_352; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_337 <= confReg_353; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_338 <= confReg_354; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_339 <= confReg_355; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_340 <= confReg_356; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_341 <= confReg_357; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_342 <= confReg_358; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_343 <= confReg_359; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_344 <= confReg_360; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_345 <= confReg_361; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_346 <= confReg_362; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_347 <= confReg_363; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_348 <= confReg_364; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_349 <= confReg_365; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_350 <= confReg_366; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_351 <= confReg_367; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_352 <= confReg_368; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_353 <= confReg_369; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_354 <= confReg_370; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_355 <= confReg_371; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_356 <= confReg_372; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_357 <= confReg_373; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_358 <= confReg_374; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_359 <= confReg_375; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_360 <= confReg_376; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_361 <= confReg_377; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_362 <= confReg_378; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_363 <= confReg_379; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_364 <= confReg_380; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_365 <= confReg_381; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_366 <= confReg_382; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_367 <= confReg_383; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_368 <= confReg_384; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_369 <= confReg_385; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_370 <= confReg_386; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_371 <= confReg_387; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_372 <= confReg_388; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_373 <= confReg_389; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_374 <= confReg_390; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_375 <= confReg_391; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_376 <= confReg_392; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_377 <= confReg_393; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_378 <= confReg_394; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_379 <= confReg_395; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_380 <= confReg_396; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_381 <= confReg_397; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_382 <= confReg_398; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_383 <= confReg_399; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_384 <= confReg_400; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_385 <= confReg_401; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_386 <= confReg_402; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_387 <= confReg_403; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_388 <= confReg_404; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_389 <= confReg_405; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_390 <= confReg_406; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_391 <= confReg_407; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_392 <= confReg_408; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_393 <= confReg_409; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_394 <= confReg_410; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_395 <= confReg_411; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_396 <= confReg_412; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_397 <= confReg_413; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_398 <= confReg_414; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_399 <= confReg_415; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_400 <= confReg_416; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_401 <= confReg_417; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_402 <= confReg_418; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_403 <= confReg_419; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_404 <= confReg_420; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_405 <= confReg_421; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_406 <= confReg_422; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_407 <= confReg_423; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_408 <= confReg_424; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_409 <= confReg_425; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_410 <= confReg_426; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_411 <= confReg_427; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_412 <= confReg_428; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_413 <= confReg_429; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_414 <= confReg_430; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_415 <= confReg_431; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_416 <= confReg_432; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_417 <= confReg_433; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_418 <= confReg_434; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_419 <= confReg_435; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_420 <= confReg_436; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_421 <= confReg_437; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_422 <= confReg_438; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_423 <= confReg_439; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_424 <= confReg_440; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_425 <= confReg_441; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_426 <= confReg_442; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_427 <= confReg_443; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_428 <= confReg_444; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_429 <= confReg_445; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_430 <= confReg_446; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_431 <= confReg_447; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_432 <= confReg_448; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_433 <= confReg_449; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_434 <= confReg_450; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_435 <= confReg_451; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_436 <= confReg_452; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_437 <= confReg_453; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_438 <= confReg_454; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_439 <= confReg_455; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_440 <= confReg_456; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_441 <= confReg_457; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_442 <= confReg_458; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_443 <= confReg_459; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_444 <= confReg_460; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_445 <= confReg_461; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_446 <= confReg_462; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_447 <= confReg_463; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_448 <= confReg_464; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_449 <= confReg_465; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_450 <= confReg_466; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_451 <= confReg_467; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_452 <= confReg_468; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_453 <= confReg_469; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_454 <= confReg_470; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_455 <= confReg_471; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_456 <= confReg_472; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_457 <= confReg_473; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_458 <= confReg_474; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_459 <= confReg_475; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_460 <= confReg_476; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_461 <= confReg_477; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_462 <= confReg_478; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_463 <= confReg_479; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_464 <= confReg_480; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_465 <= confReg_481; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_466 <= confReg_482; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_467 <= confReg_483; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_468 <= confReg_484; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_469 <= confReg_485; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_470 <= confReg_486; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_471 <= confReg_487; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_472 <= confReg_488; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_473 <= confReg_489; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_474 <= confReg_490; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_475 <= confReg_491; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_476 <= confReg_492; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_477 <= confReg_493; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_478 <= confReg_494; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_479 <= confReg_495; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_480 <= confReg_496; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_481 <= confReg_497; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_482 <= confReg_498; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_483 <= confReg_499; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_484 <= confReg_500; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_485 <= confReg_501; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_486 <= confReg_502; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_487 <= confReg_503; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_488 <= confReg_504; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_489 <= confReg_505; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_490 <= confReg_506; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_491 <= confReg_507; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_492 <= confReg_508; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_493 <= confReg_509; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_494 <= confReg_510; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_495 <= confReg_511; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_496 <= ioBundle_scan_in[0]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_497 <= ioBundle_scan_in[1]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_498 <= ioBundle_scan_in[2]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_499 <= ioBundle_scan_in[3]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_500 <= ioBundle_scan_in[4]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_501 <= ioBundle_scan_in[5]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_502 <= ioBundle_scan_in[6]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_503 <= ioBundle_scan_in[7]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_504 <= ioBundle_scan_in[8]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_505 <= ioBundle_scan_in[9]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_506 <= ioBundle_scan_in[10]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_507 <= ioBundle_scan_in[11]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_508 <= ioBundle_scan_in[12]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_509 <= ioBundle_scan_in[13]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_510 <= ioBundle_scan_in[14]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_511 <= ioBundle_scan_in[15]; // @[ScanConf.scala 38:72]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  confReg_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  confReg_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  confReg_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  confReg_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  confReg_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  confReg_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  confReg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  confReg_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  confReg_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  confReg_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  confReg_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  confReg_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  confReg_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  confReg_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  confReg_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  confReg_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  confReg_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  confReg_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  confReg_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  confReg_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  confReg_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  confReg_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  confReg_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  confReg_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  confReg_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  confReg_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  confReg_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  confReg_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  confReg_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  confReg_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  confReg_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  confReg_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  confReg_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  confReg_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  confReg_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  confReg_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  confReg_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  confReg_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  confReg_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  confReg_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  confReg_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  confReg_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  confReg_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  confReg_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  confReg_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  confReg_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  confReg_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  confReg_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  confReg_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  confReg_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  confReg_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  confReg_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  confReg_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  confReg_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  confReg_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  confReg_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  confReg_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  confReg_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  confReg_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  confReg_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  confReg_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  confReg_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  confReg_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  confReg_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  confReg_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  confReg_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  confReg_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  confReg_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  confReg_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  confReg_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  confReg_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  confReg_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  confReg_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  confReg_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  confReg_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  confReg_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  confReg_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  confReg_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  confReg_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  confReg_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  confReg_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  confReg_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  confReg_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  confReg_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  confReg_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  confReg_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  confReg_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  confReg_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  confReg_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  confReg_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  confReg_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  confReg_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  confReg_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  confReg_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  confReg_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  confReg_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  confReg_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  confReg_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  confReg_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  confReg_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  confReg_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  confReg_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  confReg_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  confReg_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  confReg_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  confReg_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  confReg_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  confReg_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  confReg_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  confReg_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  confReg_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  confReg_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  confReg_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  confReg_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  confReg_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  confReg_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  confReg_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  confReg_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  confReg_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  confReg_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  confReg_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  confReg_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  confReg_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  confReg_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  confReg_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  confReg_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  confReg_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  confReg_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  confReg_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  confReg_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  confReg_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  confReg_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  confReg_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  confReg_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  confReg_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  confReg_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  confReg_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  confReg_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  confReg_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  confReg_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  confReg_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  confReg_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  confReg_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  confReg_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  confReg_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  confReg_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  confReg_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  confReg_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  confReg_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  confReg_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  confReg_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  confReg_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  confReg_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  confReg_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  confReg_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  confReg_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  confReg_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  confReg_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  confReg_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  confReg_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  confReg_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  confReg_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  confReg_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  confReg_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  confReg_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  confReg_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  confReg_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  confReg_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  confReg_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  confReg_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  confReg_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  confReg_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  confReg_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  confReg_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  confReg_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  confReg_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  confReg_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  confReg_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  confReg_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  confReg_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  confReg_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  confReg_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  confReg_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  confReg_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  confReg_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  confReg_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  confReg_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  confReg_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  confReg_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  confReg_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  confReg_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  confReg_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  confReg_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  confReg_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  confReg_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  confReg_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  confReg_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  confReg_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  confReg_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  confReg_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  confReg_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  confReg_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  confReg_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  confReg_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  confReg_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  confReg_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  confReg_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  confReg_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  confReg_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  confReg_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  confReg_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  confReg_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  confReg_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  confReg_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  confReg_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  confReg_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  confReg_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  confReg_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  confReg_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  confReg_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  confReg_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  confReg_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  confReg_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  confReg_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  confReg_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  confReg_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  confReg_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  confReg_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  confReg_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  confReg_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  confReg_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  confReg_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  confReg_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  confReg_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  confReg_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  confReg_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  confReg_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  confReg_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  confReg_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  confReg_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  confReg_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  confReg_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  confReg_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  confReg_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  confReg_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  confReg_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  confReg_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  confReg_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  confReg_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  confReg_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  confReg_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  confReg_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  confReg_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  confReg_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  confReg_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  confReg_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  confReg_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  confReg_257 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  confReg_258 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  confReg_259 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  confReg_260 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  confReg_261 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  confReg_262 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  confReg_263 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  confReg_264 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  confReg_265 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  confReg_266 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  confReg_267 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  confReg_268 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  confReg_269 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  confReg_270 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  confReg_271 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  confReg_272 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  confReg_273 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  confReg_274 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  confReg_275 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  confReg_276 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  confReg_277 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  confReg_278 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  confReg_279 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  confReg_280 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  confReg_281 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  confReg_282 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  confReg_283 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  confReg_284 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  confReg_285 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  confReg_286 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  confReg_287 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  confReg_288 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  confReg_289 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  confReg_290 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  confReg_291 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  confReg_292 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  confReg_293 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  confReg_294 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  confReg_295 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  confReg_296 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  confReg_297 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  confReg_298 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  confReg_299 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  confReg_300 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  confReg_301 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  confReg_302 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  confReg_303 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  confReg_304 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  confReg_305 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  confReg_306 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  confReg_307 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  confReg_308 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  confReg_309 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  confReg_310 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  confReg_311 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  confReg_312 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  confReg_313 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  confReg_314 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  confReg_315 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  confReg_316 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  confReg_317 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  confReg_318 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  confReg_319 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  confReg_320 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  confReg_321 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  confReg_322 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  confReg_323 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  confReg_324 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  confReg_325 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  confReg_326 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  confReg_327 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  confReg_328 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  confReg_329 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  confReg_330 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  confReg_331 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  confReg_332 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  confReg_333 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  confReg_334 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  confReg_335 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  confReg_336 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  confReg_337 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  confReg_338 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  confReg_339 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  confReg_340 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  confReg_341 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  confReg_342 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  confReg_343 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  confReg_344 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  confReg_345 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  confReg_346 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  confReg_347 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  confReg_348 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  confReg_349 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  confReg_350 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  confReg_351 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  confReg_352 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  confReg_353 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  confReg_354 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  confReg_355 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  confReg_356 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  confReg_357 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  confReg_358 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  confReg_359 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  confReg_360 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  confReg_361 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  confReg_362 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  confReg_363 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  confReg_364 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  confReg_365 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  confReg_366 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  confReg_367 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  confReg_368 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  confReg_369 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  confReg_370 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  confReg_371 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  confReg_372 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  confReg_373 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  confReg_374 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  confReg_375 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  confReg_376 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  confReg_377 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  confReg_378 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  confReg_379 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  confReg_380 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  confReg_381 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  confReg_382 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  confReg_383 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  confReg_384 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  confReg_385 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  confReg_386 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  confReg_387 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  confReg_388 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  confReg_389 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  confReg_390 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  confReg_391 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  confReg_392 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  confReg_393 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  confReg_394 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  confReg_395 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  confReg_396 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  confReg_397 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  confReg_398 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  confReg_399 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  confReg_400 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  confReg_401 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  confReg_402 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  confReg_403 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  confReg_404 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  confReg_405 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  confReg_406 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  confReg_407 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  confReg_408 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  confReg_409 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  confReg_410 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  confReg_411 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  confReg_412 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  confReg_413 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  confReg_414 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  confReg_415 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  confReg_416 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  confReg_417 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  confReg_418 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  confReg_419 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  confReg_420 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  confReg_421 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  confReg_422 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  confReg_423 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  confReg_424 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  confReg_425 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  confReg_426 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  confReg_427 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  confReg_428 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  confReg_429 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  confReg_430 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  confReg_431 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  confReg_432 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  confReg_433 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  confReg_434 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  confReg_435 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  confReg_436 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  confReg_437 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  confReg_438 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  confReg_439 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  confReg_440 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  confReg_441 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  confReg_442 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  confReg_443 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  confReg_444 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  confReg_445 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  confReg_446 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  confReg_447 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  confReg_448 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  confReg_449 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  confReg_450 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  confReg_451 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  confReg_452 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  confReg_453 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  confReg_454 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  confReg_455 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  confReg_456 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  confReg_457 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  confReg_458 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  confReg_459 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  confReg_460 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  confReg_461 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  confReg_462 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  confReg_463 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  confReg_464 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  confReg_465 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  confReg_466 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  confReg_467 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  confReg_468 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  confReg_469 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  confReg_470 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  confReg_471 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  confReg_472 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  confReg_473 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  confReg_474 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  confReg_475 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  confReg_476 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  confReg_477 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  confReg_478 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  confReg_479 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  confReg_480 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  confReg_481 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  confReg_482 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  confReg_483 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  confReg_484 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  confReg_485 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  confReg_486 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  confReg_487 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  confReg_488 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  confReg_489 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  confReg_490 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  confReg_491 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  confReg_492 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  confReg_493 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  confReg_494 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  confReg_495 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  confReg_496 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  confReg_497 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  confReg_498 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  confReg_499 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  confReg_500 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  confReg_501 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  confReg_502 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  confReg_503 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  confReg_504 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  confReg_505 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  confReg_506 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  confReg_507 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  confReg_508 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  confReg_509 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  confReg_510 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  confReg_511 = _RAND_511[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
