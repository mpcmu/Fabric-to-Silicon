module ScanConf_Tile_11_0_EMPTY(
  input          clock,
  input          reset,
  output [287:0] ioBundle_confOut,
  input  [15:0]  ioBundle_scan_in,
  input          ioBundle_scan_en,
  output [15:0]  ioBundle_scan_out,
  input          ioBundle_scan_ioLatchEnb
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
`endif // RANDOMIZE_REG_INIT
  wire  b0mlcn000hn1n02x5_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_1_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_1_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_1_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_2_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_2_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_2_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_3_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_3_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_3_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_4_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_4_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_4_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_5_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_5_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_5_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_6_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_6_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_6_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_7_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_7_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_7_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_8_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_8_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_8_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_9_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_9_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_9_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_10_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_10_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_10_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_11_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_11_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_11_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_12_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_12_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_12_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_13_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_13_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_13_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_14_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_14_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_14_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_15_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_15_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_15_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_16_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_16_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_16_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_17_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_17_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_17_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_18_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_18_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_18_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_19_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_19_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_19_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_20_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_20_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_20_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_21_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_21_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_21_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_22_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_22_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_22_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_23_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_23_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_23_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_24_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_24_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_24_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_25_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_25_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_25_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_26_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_26_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_26_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_27_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_27_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_27_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_28_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_28_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_28_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_29_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_29_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_29_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_30_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_30_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_30_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_31_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_31_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_31_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_32_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_32_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_32_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_33_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_33_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_33_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_34_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_34_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_34_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_35_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_35_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_35_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_36_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_36_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_36_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_37_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_37_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_37_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_38_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_38_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_38_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_39_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_39_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_39_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_40_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_40_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_40_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_41_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_41_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_41_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_42_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_42_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_42_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_43_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_43_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_43_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_44_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_44_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_44_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_45_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_45_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_45_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_46_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_46_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_46_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_47_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_47_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_47_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_48_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_48_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_48_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_49_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_49_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_49_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_50_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_50_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_50_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_51_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_51_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_51_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_52_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_52_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_52_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_53_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_53_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_53_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_54_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_54_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_54_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_55_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_55_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_55_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_56_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_56_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_56_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_57_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_57_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_57_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_58_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_58_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_58_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_59_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_59_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_59_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_60_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_60_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_60_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_61_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_61_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_61_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_62_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_62_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_62_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_63_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_63_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_63_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_64_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_64_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_64_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_65_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_65_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_65_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_66_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_66_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_66_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_67_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_67_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_67_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_68_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_68_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_68_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_69_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_69_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_69_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_70_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_70_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_70_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_71_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_71_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_71_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_72_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_72_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_72_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_73_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_73_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_73_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_74_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_74_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_74_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_75_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_75_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_75_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_76_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_76_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_76_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_77_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_77_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_77_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_78_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_78_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_78_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_79_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_79_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_79_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_80_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_80_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_80_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_81_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_81_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_81_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_82_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_82_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_82_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_83_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_83_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_83_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_84_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_84_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_84_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_85_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_85_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_85_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_86_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_86_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_86_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_87_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_87_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_87_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_88_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_88_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_88_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_89_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_89_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_89_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_90_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_90_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_90_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_91_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_91_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_91_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_92_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_92_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_92_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_93_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_93_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_93_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_94_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_94_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_94_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_95_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_95_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_95_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_96_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_96_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_96_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_97_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_97_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_97_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_98_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_98_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_98_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_99_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_99_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_99_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_100_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_100_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_100_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_101_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_101_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_101_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_102_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_102_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_102_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_103_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_103_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_103_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_104_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_104_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_104_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_105_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_105_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_105_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_106_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_106_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_106_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_107_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_107_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_107_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_108_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_108_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_108_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_109_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_109_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_109_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_110_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_110_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_110_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_111_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_111_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_111_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_112_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_112_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_112_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_113_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_113_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_113_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_114_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_114_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_114_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_115_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_115_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_115_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_116_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_116_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_116_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_117_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_117_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_117_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_118_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_118_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_118_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_119_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_119_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_119_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_120_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_120_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_120_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_121_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_121_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_121_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_122_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_122_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_122_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_123_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_123_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_123_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_124_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_124_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_124_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_125_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_125_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_125_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_126_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_126_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_126_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_127_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_127_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_127_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_128_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_128_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_128_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_129_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_129_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_129_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_130_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_130_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_130_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_131_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_131_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_131_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_132_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_132_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_132_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_133_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_133_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_133_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_134_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_134_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_134_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_135_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_135_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_135_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_136_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_136_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_136_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_137_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_137_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_137_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_138_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_138_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_138_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_139_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_139_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_139_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_140_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_140_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_140_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_141_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_141_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_141_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_142_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_142_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_142_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_143_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_143_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_143_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_144_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_144_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_144_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_145_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_145_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_145_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_146_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_146_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_146_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_147_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_147_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_147_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_148_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_148_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_148_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_149_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_149_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_149_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_150_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_150_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_150_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_151_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_151_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_151_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_152_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_152_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_152_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_153_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_153_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_153_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_154_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_154_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_154_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_155_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_155_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_155_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_156_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_156_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_156_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_157_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_157_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_157_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_158_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_158_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_158_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_159_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_159_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_159_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_160_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_160_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_160_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_161_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_161_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_161_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_162_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_162_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_162_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_163_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_163_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_163_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_164_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_164_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_164_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_165_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_165_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_165_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_166_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_166_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_166_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_167_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_167_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_167_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_168_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_168_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_168_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_169_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_169_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_169_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_170_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_170_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_170_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_171_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_171_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_171_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_172_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_172_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_172_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_173_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_173_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_173_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_174_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_174_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_174_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_175_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_175_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_175_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_176_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_176_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_176_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_177_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_177_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_177_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_178_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_178_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_178_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_179_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_179_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_179_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_180_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_180_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_180_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_181_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_181_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_181_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_182_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_182_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_182_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_183_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_183_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_183_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_184_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_184_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_184_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_185_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_185_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_185_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_186_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_186_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_186_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_187_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_187_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_187_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_188_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_188_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_188_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_189_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_189_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_189_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_190_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_190_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_190_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_191_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_191_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_191_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_192_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_192_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_192_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_193_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_193_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_193_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_194_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_194_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_194_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_195_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_195_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_195_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_196_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_196_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_196_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_197_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_197_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_197_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_198_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_198_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_198_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_199_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_199_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_199_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_200_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_200_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_200_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_201_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_201_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_201_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_202_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_202_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_202_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_203_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_203_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_203_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_204_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_204_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_204_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_205_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_205_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_205_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_206_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_206_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_206_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_207_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_207_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_207_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_208_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_208_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_208_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_209_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_209_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_209_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_210_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_210_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_210_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_211_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_211_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_211_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_212_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_212_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_212_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_213_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_213_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_213_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_214_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_214_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_214_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_215_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_215_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_215_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_216_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_216_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_216_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_217_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_217_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_217_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_218_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_218_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_218_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_219_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_219_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_219_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_220_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_220_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_220_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_221_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_221_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_221_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_222_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_222_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_222_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_223_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_223_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_223_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_224_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_224_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_224_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_225_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_225_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_225_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_226_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_226_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_226_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_227_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_227_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_227_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_228_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_228_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_228_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_229_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_229_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_229_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_230_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_230_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_230_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_231_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_231_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_231_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_232_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_232_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_232_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_233_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_233_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_233_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_234_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_234_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_234_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_235_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_235_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_235_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_236_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_236_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_236_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_237_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_237_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_237_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_238_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_238_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_238_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_239_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_239_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_239_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_240_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_240_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_240_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_241_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_241_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_241_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_242_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_242_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_242_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_243_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_243_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_243_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_244_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_244_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_244_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_245_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_245_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_245_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_246_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_246_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_246_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_247_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_247_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_247_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_248_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_248_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_248_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_249_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_249_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_249_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_250_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_250_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_250_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_251_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_251_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_251_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_252_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_252_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_252_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_253_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_253_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_253_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_254_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_254_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_254_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_255_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_255_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_255_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_256_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_256_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_256_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_257_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_257_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_257_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_258_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_258_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_258_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_259_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_259_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_259_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_260_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_260_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_260_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_261_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_261_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_261_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_262_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_262_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_262_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_263_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_263_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_263_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_264_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_264_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_264_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_265_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_265_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_265_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_266_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_266_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_266_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_267_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_267_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_267_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_268_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_268_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_268_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_269_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_269_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_269_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_270_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_270_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_270_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_271_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_271_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_271_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_272_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_272_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_272_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_273_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_273_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_273_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_274_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_274_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_274_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_275_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_275_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_275_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_276_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_276_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_276_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_277_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_277_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_277_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_278_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_278_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_278_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_279_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_279_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_279_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_280_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_280_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_280_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_281_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_281_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_281_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_282_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_282_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_282_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_283_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_283_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_283_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_284_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_284_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_284_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_285_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_285_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_285_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_286_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_286_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_286_o; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_287_d; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_287_clk; // @[ScanConfRadh.scala 61:46]
  wire  b0mlcn000hn1n02x5_287_o; // @[ScanConfRadh.scala 61:46]
  reg  confReg_0; // @[ScanConfRadh.scala 45:20]
  reg  confReg_1; // @[ScanConfRadh.scala 45:20]
  reg  confReg_2; // @[ScanConfRadh.scala 45:20]
  reg  confReg_3; // @[ScanConfRadh.scala 45:20]
  reg  confReg_4; // @[ScanConfRadh.scala 45:20]
  reg  confReg_5; // @[ScanConfRadh.scala 45:20]
  reg  confReg_6; // @[ScanConfRadh.scala 45:20]
  reg  confReg_7; // @[ScanConfRadh.scala 45:20]
  reg  confReg_8; // @[ScanConfRadh.scala 45:20]
  reg  confReg_9; // @[ScanConfRadh.scala 45:20]
  reg  confReg_10; // @[ScanConfRadh.scala 45:20]
  reg  confReg_11; // @[ScanConfRadh.scala 45:20]
  reg  confReg_12; // @[ScanConfRadh.scala 45:20]
  reg  confReg_13; // @[ScanConfRadh.scala 45:20]
  reg  confReg_14; // @[ScanConfRadh.scala 45:20]
  reg  confReg_15; // @[ScanConfRadh.scala 45:20]
  reg  confReg_16; // @[ScanConfRadh.scala 45:20]
  reg  confReg_17; // @[ScanConfRadh.scala 45:20]
  reg  confReg_18; // @[ScanConfRadh.scala 45:20]
  reg  confReg_19; // @[ScanConfRadh.scala 45:20]
  reg  confReg_20; // @[ScanConfRadh.scala 45:20]
  reg  confReg_21; // @[ScanConfRadh.scala 45:20]
  reg  confReg_22; // @[ScanConfRadh.scala 45:20]
  reg  confReg_23; // @[ScanConfRadh.scala 45:20]
  reg  confReg_24; // @[ScanConfRadh.scala 45:20]
  reg  confReg_25; // @[ScanConfRadh.scala 45:20]
  reg  confReg_26; // @[ScanConfRadh.scala 45:20]
  reg  confReg_27; // @[ScanConfRadh.scala 45:20]
  reg  confReg_28; // @[ScanConfRadh.scala 45:20]
  reg  confReg_29; // @[ScanConfRadh.scala 45:20]
  reg  confReg_30; // @[ScanConfRadh.scala 45:20]
  reg  confReg_31; // @[ScanConfRadh.scala 45:20]
  reg  confReg_32; // @[ScanConfRadh.scala 45:20]
  reg  confReg_33; // @[ScanConfRadh.scala 45:20]
  reg  confReg_34; // @[ScanConfRadh.scala 45:20]
  reg  confReg_35; // @[ScanConfRadh.scala 45:20]
  reg  confReg_36; // @[ScanConfRadh.scala 45:20]
  reg  confReg_37; // @[ScanConfRadh.scala 45:20]
  reg  confReg_38; // @[ScanConfRadh.scala 45:20]
  reg  confReg_39; // @[ScanConfRadh.scala 45:20]
  reg  confReg_40; // @[ScanConfRadh.scala 45:20]
  reg  confReg_41; // @[ScanConfRadh.scala 45:20]
  reg  confReg_42; // @[ScanConfRadh.scala 45:20]
  reg  confReg_43; // @[ScanConfRadh.scala 45:20]
  reg  confReg_44; // @[ScanConfRadh.scala 45:20]
  reg  confReg_45; // @[ScanConfRadh.scala 45:20]
  reg  confReg_46; // @[ScanConfRadh.scala 45:20]
  reg  confReg_47; // @[ScanConfRadh.scala 45:20]
  reg  confReg_48; // @[ScanConfRadh.scala 45:20]
  reg  confReg_49; // @[ScanConfRadh.scala 45:20]
  reg  confReg_50; // @[ScanConfRadh.scala 45:20]
  reg  confReg_51; // @[ScanConfRadh.scala 45:20]
  reg  confReg_52; // @[ScanConfRadh.scala 45:20]
  reg  confReg_53; // @[ScanConfRadh.scala 45:20]
  reg  confReg_54; // @[ScanConfRadh.scala 45:20]
  reg  confReg_55; // @[ScanConfRadh.scala 45:20]
  reg  confReg_56; // @[ScanConfRadh.scala 45:20]
  reg  confReg_57; // @[ScanConfRadh.scala 45:20]
  reg  confReg_58; // @[ScanConfRadh.scala 45:20]
  reg  confReg_59; // @[ScanConfRadh.scala 45:20]
  reg  confReg_60; // @[ScanConfRadh.scala 45:20]
  reg  confReg_61; // @[ScanConfRadh.scala 45:20]
  reg  confReg_62; // @[ScanConfRadh.scala 45:20]
  reg  confReg_63; // @[ScanConfRadh.scala 45:20]
  reg  confReg_64; // @[ScanConfRadh.scala 45:20]
  reg  confReg_65; // @[ScanConfRadh.scala 45:20]
  reg  confReg_66; // @[ScanConfRadh.scala 45:20]
  reg  confReg_67; // @[ScanConfRadh.scala 45:20]
  reg  confReg_68; // @[ScanConfRadh.scala 45:20]
  reg  confReg_69; // @[ScanConfRadh.scala 45:20]
  reg  confReg_70; // @[ScanConfRadh.scala 45:20]
  reg  confReg_71; // @[ScanConfRadh.scala 45:20]
  reg  confReg_72; // @[ScanConfRadh.scala 45:20]
  reg  confReg_73; // @[ScanConfRadh.scala 45:20]
  reg  confReg_74; // @[ScanConfRadh.scala 45:20]
  reg  confReg_75; // @[ScanConfRadh.scala 45:20]
  reg  confReg_76; // @[ScanConfRadh.scala 45:20]
  reg  confReg_77; // @[ScanConfRadh.scala 45:20]
  reg  confReg_78; // @[ScanConfRadh.scala 45:20]
  reg  confReg_79; // @[ScanConfRadh.scala 45:20]
  reg  confReg_80; // @[ScanConfRadh.scala 45:20]
  reg  confReg_81; // @[ScanConfRadh.scala 45:20]
  reg  confReg_82; // @[ScanConfRadh.scala 45:20]
  reg  confReg_83; // @[ScanConfRadh.scala 45:20]
  reg  confReg_84; // @[ScanConfRadh.scala 45:20]
  reg  confReg_85; // @[ScanConfRadh.scala 45:20]
  reg  confReg_86; // @[ScanConfRadh.scala 45:20]
  reg  confReg_87; // @[ScanConfRadh.scala 45:20]
  reg  confReg_88; // @[ScanConfRadh.scala 45:20]
  reg  confReg_89; // @[ScanConfRadh.scala 45:20]
  reg  confReg_90; // @[ScanConfRadh.scala 45:20]
  reg  confReg_91; // @[ScanConfRadh.scala 45:20]
  reg  confReg_92; // @[ScanConfRadh.scala 45:20]
  reg  confReg_93; // @[ScanConfRadh.scala 45:20]
  reg  confReg_94; // @[ScanConfRadh.scala 45:20]
  reg  confReg_95; // @[ScanConfRadh.scala 45:20]
  reg  confReg_96; // @[ScanConfRadh.scala 45:20]
  reg  confReg_97; // @[ScanConfRadh.scala 45:20]
  reg  confReg_98; // @[ScanConfRadh.scala 45:20]
  reg  confReg_99; // @[ScanConfRadh.scala 45:20]
  reg  confReg_100; // @[ScanConfRadh.scala 45:20]
  reg  confReg_101; // @[ScanConfRadh.scala 45:20]
  reg  confReg_102; // @[ScanConfRadh.scala 45:20]
  reg  confReg_103; // @[ScanConfRadh.scala 45:20]
  reg  confReg_104; // @[ScanConfRadh.scala 45:20]
  reg  confReg_105; // @[ScanConfRadh.scala 45:20]
  reg  confReg_106; // @[ScanConfRadh.scala 45:20]
  reg  confReg_107; // @[ScanConfRadh.scala 45:20]
  reg  confReg_108; // @[ScanConfRadh.scala 45:20]
  reg  confReg_109; // @[ScanConfRadh.scala 45:20]
  reg  confReg_110; // @[ScanConfRadh.scala 45:20]
  reg  confReg_111; // @[ScanConfRadh.scala 45:20]
  reg  confReg_112; // @[ScanConfRadh.scala 45:20]
  reg  confReg_113; // @[ScanConfRadh.scala 45:20]
  reg  confReg_114; // @[ScanConfRadh.scala 45:20]
  reg  confReg_115; // @[ScanConfRadh.scala 45:20]
  reg  confReg_116; // @[ScanConfRadh.scala 45:20]
  reg  confReg_117; // @[ScanConfRadh.scala 45:20]
  reg  confReg_118; // @[ScanConfRadh.scala 45:20]
  reg  confReg_119; // @[ScanConfRadh.scala 45:20]
  reg  confReg_120; // @[ScanConfRadh.scala 45:20]
  reg  confReg_121; // @[ScanConfRadh.scala 45:20]
  reg  confReg_122; // @[ScanConfRadh.scala 45:20]
  reg  confReg_123; // @[ScanConfRadh.scala 45:20]
  reg  confReg_124; // @[ScanConfRadh.scala 45:20]
  reg  confReg_125; // @[ScanConfRadh.scala 45:20]
  reg  confReg_126; // @[ScanConfRadh.scala 45:20]
  reg  confReg_127; // @[ScanConfRadh.scala 45:20]
  reg  confReg_128; // @[ScanConfRadh.scala 45:20]
  reg  confReg_129; // @[ScanConfRadh.scala 45:20]
  reg  confReg_130; // @[ScanConfRadh.scala 45:20]
  reg  confReg_131; // @[ScanConfRadh.scala 45:20]
  reg  confReg_132; // @[ScanConfRadh.scala 45:20]
  reg  confReg_133; // @[ScanConfRadh.scala 45:20]
  reg  confReg_134; // @[ScanConfRadh.scala 45:20]
  reg  confReg_135; // @[ScanConfRadh.scala 45:20]
  reg  confReg_136; // @[ScanConfRadh.scala 45:20]
  reg  confReg_137; // @[ScanConfRadh.scala 45:20]
  reg  confReg_138; // @[ScanConfRadh.scala 45:20]
  reg  confReg_139; // @[ScanConfRadh.scala 45:20]
  reg  confReg_140; // @[ScanConfRadh.scala 45:20]
  reg  confReg_141; // @[ScanConfRadh.scala 45:20]
  reg  confReg_142; // @[ScanConfRadh.scala 45:20]
  reg  confReg_143; // @[ScanConfRadh.scala 45:20]
  reg  confReg_144; // @[ScanConfRadh.scala 45:20]
  reg  confReg_145; // @[ScanConfRadh.scala 45:20]
  reg  confReg_146; // @[ScanConfRadh.scala 45:20]
  reg  confReg_147; // @[ScanConfRadh.scala 45:20]
  reg  confReg_148; // @[ScanConfRadh.scala 45:20]
  reg  confReg_149; // @[ScanConfRadh.scala 45:20]
  reg  confReg_150; // @[ScanConfRadh.scala 45:20]
  reg  confReg_151; // @[ScanConfRadh.scala 45:20]
  reg  confReg_152; // @[ScanConfRadh.scala 45:20]
  reg  confReg_153; // @[ScanConfRadh.scala 45:20]
  reg  confReg_154; // @[ScanConfRadh.scala 45:20]
  reg  confReg_155; // @[ScanConfRadh.scala 45:20]
  reg  confReg_156; // @[ScanConfRadh.scala 45:20]
  reg  confReg_157; // @[ScanConfRadh.scala 45:20]
  reg  confReg_158; // @[ScanConfRadh.scala 45:20]
  reg  confReg_159; // @[ScanConfRadh.scala 45:20]
  reg  confReg_160; // @[ScanConfRadh.scala 45:20]
  reg  confReg_161; // @[ScanConfRadh.scala 45:20]
  reg  confReg_162; // @[ScanConfRadh.scala 45:20]
  reg  confReg_163; // @[ScanConfRadh.scala 45:20]
  reg  confReg_164; // @[ScanConfRadh.scala 45:20]
  reg  confReg_165; // @[ScanConfRadh.scala 45:20]
  reg  confReg_166; // @[ScanConfRadh.scala 45:20]
  reg  confReg_167; // @[ScanConfRadh.scala 45:20]
  reg  confReg_168; // @[ScanConfRadh.scala 45:20]
  reg  confReg_169; // @[ScanConfRadh.scala 45:20]
  reg  confReg_170; // @[ScanConfRadh.scala 45:20]
  reg  confReg_171; // @[ScanConfRadh.scala 45:20]
  reg  confReg_172; // @[ScanConfRadh.scala 45:20]
  reg  confReg_173; // @[ScanConfRadh.scala 45:20]
  reg  confReg_174; // @[ScanConfRadh.scala 45:20]
  reg  confReg_175; // @[ScanConfRadh.scala 45:20]
  reg  confReg_176; // @[ScanConfRadh.scala 45:20]
  reg  confReg_177; // @[ScanConfRadh.scala 45:20]
  reg  confReg_178; // @[ScanConfRadh.scala 45:20]
  reg  confReg_179; // @[ScanConfRadh.scala 45:20]
  reg  confReg_180; // @[ScanConfRadh.scala 45:20]
  reg  confReg_181; // @[ScanConfRadh.scala 45:20]
  reg  confReg_182; // @[ScanConfRadh.scala 45:20]
  reg  confReg_183; // @[ScanConfRadh.scala 45:20]
  reg  confReg_184; // @[ScanConfRadh.scala 45:20]
  reg  confReg_185; // @[ScanConfRadh.scala 45:20]
  reg  confReg_186; // @[ScanConfRadh.scala 45:20]
  reg  confReg_187; // @[ScanConfRadh.scala 45:20]
  reg  confReg_188; // @[ScanConfRadh.scala 45:20]
  reg  confReg_189; // @[ScanConfRadh.scala 45:20]
  reg  confReg_190; // @[ScanConfRadh.scala 45:20]
  reg  confReg_191; // @[ScanConfRadh.scala 45:20]
  reg  confReg_192; // @[ScanConfRadh.scala 45:20]
  reg  confReg_193; // @[ScanConfRadh.scala 45:20]
  reg  confReg_194; // @[ScanConfRadh.scala 45:20]
  reg  confReg_195; // @[ScanConfRadh.scala 45:20]
  reg  confReg_196; // @[ScanConfRadh.scala 45:20]
  reg  confReg_197; // @[ScanConfRadh.scala 45:20]
  reg  confReg_198; // @[ScanConfRadh.scala 45:20]
  reg  confReg_199; // @[ScanConfRadh.scala 45:20]
  reg  confReg_200; // @[ScanConfRadh.scala 45:20]
  reg  confReg_201; // @[ScanConfRadh.scala 45:20]
  reg  confReg_202; // @[ScanConfRadh.scala 45:20]
  reg  confReg_203; // @[ScanConfRadh.scala 45:20]
  reg  confReg_204; // @[ScanConfRadh.scala 45:20]
  reg  confReg_205; // @[ScanConfRadh.scala 45:20]
  reg  confReg_206; // @[ScanConfRadh.scala 45:20]
  reg  confReg_207; // @[ScanConfRadh.scala 45:20]
  reg  confReg_208; // @[ScanConfRadh.scala 45:20]
  reg  confReg_209; // @[ScanConfRadh.scala 45:20]
  reg  confReg_210; // @[ScanConfRadh.scala 45:20]
  reg  confReg_211; // @[ScanConfRadh.scala 45:20]
  reg  confReg_212; // @[ScanConfRadh.scala 45:20]
  reg  confReg_213; // @[ScanConfRadh.scala 45:20]
  reg  confReg_214; // @[ScanConfRadh.scala 45:20]
  reg  confReg_215; // @[ScanConfRadh.scala 45:20]
  reg  confReg_216; // @[ScanConfRadh.scala 45:20]
  reg  confReg_217; // @[ScanConfRadh.scala 45:20]
  reg  confReg_218; // @[ScanConfRadh.scala 45:20]
  reg  confReg_219; // @[ScanConfRadh.scala 45:20]
  reg  confReg_220; // @[ScanConfRadh.scala 45:20]
  reg  confReg_221; // @[ScanConfRadh.scala 45:20]
  reg  confReg_222; // @[ScanConfRadh.scala 45:20]
  reg  confReg_223; // @[ScanConfRadh.scala 45:20]
  reg  confReg_224; // @[ScanConfRadh.scala 45:20]
  reg  confReg_225; // @[ScanConfRadh.scala 45:20]
  reg  confReg_226; // @[ScanConfRadh.scala 45:20]
  reg  confReg_227; // @[ScanConfRadh.scala 45:20]
  reg  confReg_228; // @[ScanConfRadh.scala 45:20]
  reg  confReg_229; // @[ScanConfRadh.scala 45:20]
  reg  confReg_230; // @[ScanConfRadh.scala 45:20]
  reg  confReg_231; // @[ScanConfRadh.scala 45:20]
  reg  confReg_232; // @[ScanConfRadh.scala 45:20]
  reg  confReg_233; // @[ScanConfRadh.scala 45:20]
  reg  confReg_234; // @[ScanConfRadh.scala 45:20]
  reg  confReg_235; // @[ScanConfRadh.scala 45:20]
  reg  confReg_236; // @[ScanConfRadh.scala 45:20]
  reg  confReg_237; // @[ScanConfRadh.scala 45:20]
  reg  confReg_238; // @[ScanConfRadh.scala 45:20]
  reg  confReg_239; // @[ScanConfRadh.scala 45:20]
  reg  confReg_240; // @[ScanConfRadh.scala 45:20]
  reg  confReg_241; // @[ScanConfRadh.scala 45:20]
  reg  confReg_242; // @[ScanConfRadh.scala 45:20]
  reg  confReg_243; // @[ScanConfRadh.scala 45:20]
  reg  confReg_244; // @[ScanConfRadh.scala 45:20]
  reg  confReg_245; // @[ScanConfRadh.scala 45:20]
  reg  confReg_246; // @[ScanConfRadh.scala 45:20]
  reg  confReg_247; // @[ScanConfRadh.scala 45:20]
  reg  confReg_248; // @[ScanConfRadh.scala 45:20]
  reg  confReg_249; // @[ScanConfRadh.scala 45:20]
  reg  confReg_250; // @[ScanConfRadh.scala 45:20]
  reg  confReg_251; // @[ScanConfRadh.scala 45:20]
  reg  confReg_252; // @[ScanConfRadh.scala 45:20]
  reg  confReg_253; // @[ScanConfRadh.scala 45:20]
  reg  confReg_254; // @[ScanConfRadh.scala 45:20]
  reg  confReg_255; // @[ScanConfRadh.scala 45:20]
  reg  confReg_256; // @[ScanConfRadh.scala 45:20]
  reg  confReg_257; // @[ScanConfRadh.scala 45:20]
  reg  confReg_258; // @[ScanConfRadh.scala 45:20]
  reg  confReg_259; // @[ScanConfRadh.scala 45:20]
  reg  confReg_260; // @[ScanConfRadh.scala 45:20]
  reg  confReg_261; // @[ScanConfRadh.scala 45:20]
  reg  confReg_262; // @[ScanConfRadh.scala 45:20]
  reg  confReg_263; // @[ScanConfRadh.scala 45:20]
  reg  confReg_264; // @[ScanConfRadh.scala 45:20]
  reg  confReg_265; // @[ScanConfRadh.scala 45:20]
  reg  confReg_266; // @[ScanConfRadh.scala 45:20]
  reg  confReg_267; // @[ScanConfRadh.scala 45:20]
  reg  confReg_268; // @[ScanConfRadh.scala 45:20]
  reg  confReg_269; // @[ScanConfRadh.scala 45:20]
  reg  confReg_270; // @[ScanConfRadh.scala 45:20]
  reg  confReg_271; // @[ScanConfRadh.scala 45:20]
  reg  confReg_272; // @[ScanConfRadh.scala 45:20]
  reg  confReg_273; // @[ScanConfRadh.scala 45:20]
  reg  confReg_274; // @[ScanConfRadh.scala 45:20]
  reg  confReg_275; // @[ScanConfRadh.scala 45:20]
  reg  confReg_276; // @[ScanConfRadh.scala 45:20]
  reg  confReg_277; // @[ScanConfRadh.scala 45:20]
  reg  confReg_278; // @[ScanConfRadh.scala 45:20]
  reg  confReg_279; // @[ScanConfRadh.scala 45:20]
  reg  confReg_280; // @[ScanConfRadh.scala 45:20]
  reg  confReg_281; // @[ScanConfRadh.scala 45:20]
  reg  confReg_282; // @[ScanConfRadh.scala 45:20]
  reg  confReg_283; // @[ScanConfRadh.scala 45:20]
  reg  confReg_284; // @[ScanConfRadh.scala 45:20]
  reg  confReg_285; // @[ScanConfRadh.scala 45:20]
  reg  confReg_286; // @[ScanConfRadh.scala 45:20]
  reg  confReg_287; // @[ScanConfRadh.scala 45:20]
  wire [15:0] io_scan_in = ioBundle_scan_in; // @[ScanConfRadh.scala 40:16 70:12]
  wire  _confReg_272_T = ioBundle_scan_in[0]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_273_T = ioBundle_scan_in[1]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_274_T = ioBundle_scan_in[2]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_275_T = ioBundle_scan_in[3]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_276_T = ioBundle_scan_in[4]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_277_T = ioBundle_scan_in[5]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_278_T = ioBundle_scan_in[6]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_279_T = ioBundle_scan_in[7]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_280_T = ioBundle_scan_in[8]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_281_T = ioBundle_scan_in[9]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_282_T = ioBundle_scan_in[10]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_283_T = ioBundle_scan_in[11]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_284_T = ioBundle_scan_in[12]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_285_T = ioBundle_scan_in[13]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_286_T = ioBundle_scan_in[14]; // @[ScanConfRadh.scala 51:85]
  wire  _confReg_287_T = ioBundle_scan_in[15]; // @[ScanConfRadh.scala 51:85]
  wire  io_scan_en = ioBundle_scan_en; // @[ScanConfRadh.scala 40:16 70:12]
  wire  _GEN_0 = ioBundle_scan_en ? ioBundle_scan_in[0] : confReg_272; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_1 = ioBundle_scan_en ? ioBundle_scan_in[1] : confReg_273; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_2 = ioBundle_scan_en ? ioBundle_scan_in[2] : confReg_274; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_3 = ioBundle_scan_en ? ioBundle_scan_in[3] : confReg_275; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_4 = ioBundle_scan_en ? ioBundle_scan_in[4] : confReg_276; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_5 = ioBundle_scan_en ? ioBundle_scan_in[5] : confReg_277; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_6 = ioBundle_scan_en ? ioBundle_scan_in[6] : confReg_278; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_7 = ioBundle_scan_en ? ioBundle_scan_in[7] : confReg_279; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_8 = ioBundle_scan_en ? ioBundle_scan_in[8] : confReg_280; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_9 = ioBundle_scan_en ? ioBundle_scan_in[9] : confReg_281; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_10 = ioBundle_scan_en ? ioBundle_scan_in[10] : confReg_282; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_11 = ioBundle_scan_en ? ioBundle_scan_in[11] : confReg_283; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_12 = ioBundle_scan_en ? ioBundle_scan_in[12] : confReg_284; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_13 = ioBundle_scan_en ? ioBundle_scan_in[13] : confReg_285; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_14 = ioBundle_scan_en ? ioBundle_scan_in[14] : confReg_286; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_15 = ioBundle_scan_en ? ioBundle_scan_in[15] : confReg_287; // @[ScanConfRadh.scala 45:20 50:20 51:72]
  wire  _GEN_16 = ioBundle_scan_en ? confReg_16 : confReg_0; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_17 = ioBundle_scan_en ? confReg_17 : confReg_1; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_18 = ioBundle_scan_en ? confReg_18 : confReg_2; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_19 = ioBundle_scan_en ? confReg_19 : confReg_3; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_20 = ioBundle_scan_en ? confReg_20 : confReg_4; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_21 = ioBundle_scan_en ? confReg_21 : confReg_5; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_22 = ioBundle_scan_en ? confReg_22 : confReg_6; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_23 = ioBundle_scan_en ? confReg_23 : confReg_7; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_24 = ioBundle_scan_en ? confReg_24 : confReg_8; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_25 = ioBundle_scan_en ? confReg_25 : confReg_9; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_26 = ioBundle_scan_en ? confReg_26 : confReg_10; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_27 = ioBundle_scan_en ? confReg_27 : confReg_11; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_28 = ioBundle_scan_en ? confReg_28 : confReg_12; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_29 = ioBundle_scan_en ? confReg_29 : confReg_13; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_30 = ioBundle_scan_en ? confReg_30 : confReg_14; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_31 = ioBundle_scan_en ? confReg_31 : confReg_15; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_32 = ioBundle_scan_en ? confReg_32 : confReg_16; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_33 = ioBundle_scan_en ? confReg_33 : confReg_17; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_34 = ioBundle_scan_en ? confReg_34 : confReg_18; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_35 = ioBundle_scan_en ? confReg_35 : confReg_19; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_36 = ioBundle_scan_en ? confReg_36 : confReg_20; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_37 = ioBundle_scan_en ? confReg_37 : confReg_21; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_38 = ioBundle_scan_en ? confReg_38 : confReg_22; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_39 = ioBundle_scan_en ? confReg_39 : confReg_23; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_40 = ioBundle_scan_en ? confReg_40 : confReg_24; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_41 = ioBundle_scan_en ? confReg_41 : confReg_25; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_42 = ioBundle_scan_en ? confReg_42 : confReg_26; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_43 = ioBundle_scan_en ? confReg_43 : confReg_27; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_44 = ioBundle_scan_en ? confReg_44 : confReg_28; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_45 = ioBundle_scan_en ? confReg_45 : confReg_29; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_46 = ioBundle_scan_en ? confReg_46 : confReg_30; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_47 = ioBundle_scan_en ? confReg_47 : confReg_31; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_48 = ioBundle_scan_en ? confReg_48 : confReg_32; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_49 = ioBundle_scan_en ? confReg_49 : confReg_33; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_50 = ioBundle_scan_en ? confReg_50 : confReg_34; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_51 = ioBundle_scan_en ? confReg_51 : confReg_35; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_52 = ioBundle_scan_en ? confReg_52 : confReg_36; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_53 = ioBundle_scan_en ? confReg_53 : confReg_37; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_54 = ioBundle_scan_en ? confReg_54 : confReg_38; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_55 = ioBundle_scan_en ? confReg_55 : confReg_39; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_56 = ioBundle_scan_en ? confReg_56 : confReg_40; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_57 = ioBundle_scan_en ? confReg_57 : confReg_41; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_58 = ioBundle_scan_en ? confReg_58 : confReg_42; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_59 = ioBundle_scan_en ? confReg_59 : confReg_43; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_60 = ioBundle_scan_en ? confReg_60 : confReg_44; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_61 = ioBundle_scan_en ? confReg_61 : confReg_45; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_62 = ioBundle_scan_en ? confReg_62 : confReg_46; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_63 = ioBundle_scan_en ? confReg_63 : confReg_47; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_64 = ioBundle_scan_en ? confReg_64 : confReg_48; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_65 = ioBundle_scan_en ? confReg_65 : confReg_49; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_66 = ioBundle_scan_en ? confReg_66 : confReg_50; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_67 = ioBundle_scan_en ? confReg_67 : confReg_51; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_68 = ioBundle_scan_en ? confReg_68 : confReg_52; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_69 = ioBundle_scan_en ? confReg_69 : confReg_53; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_70 = ioBundle_scan_en ? confReg_70 : confReg_54; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_71 = ioBundle_scan_en ? confReg_71 : confReg_55; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_72 = ioBundle_scan_en ? confReg_72 : confReg_56; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_73 = ioBundle_scan_en ? confReg_73 : confReg_57; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_74 = ioBundle_scan_en ? confReg_74 : confReg_58; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_75 = ioBundle_scan_en ? confReg_75 : confReg_59; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_76 = ioBundle_scan_en ? confReg_76 : confReg_60; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_77 = ioBundle_scan_en ? confReg_77 : confReg_61; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_78 = ioBundle_scan_en ? confReg_78 : confReg_62; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_79 = ioBundle_scan_en ? confReg_79 : confReg_63; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_80 = ioBundle_scan_en ? confReg_80 : confReg_64; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_81 = ioBundle_scan_en ? confReg_81 : confReg_65; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_82 = ioBundle_scan_en ? confReg_82 : confReg_66; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_83 = ioBundle_scan_en ? confReg_83 : confReg_67; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_84 = ioBundle_scan_en ? confReg_84 : confReg_68; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_85 = ioBundle_scan_en ? confReg_85 : confReg_69; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_86 = ioBundle_scan_en ? confReg_86 : confReg_70; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_87 = ioBundle_scan_en ? confReg_87 : confReg_71; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_88 = ioBundle_scan_en ? confReg_88 : confReg_72; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_89 = ioBundle_scan_en ? confReg_89 : confReg_73; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_90 = ioBundle_scan_en ? confReg_90 : confReg_74; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_91 = ioBundle_scan_en ? confReg_91 : confReg_75; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_92 = ioBundle_scan_en ? confReg_92 : confReg_76; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_93 = ioBundle_scan_en ? confReg_93 : confReg_77; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_94 = ioBundle_scan_en ? confReg_94 : confReg_78; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_95 = ioBundle_scan_en ? confReg_95 : confReg_79; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_96 = ioBundle_scan_en ? confReg_96 : confReg_80; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_97 = ioBundle_scan_en ? confReg_97 : confReg_81; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_98 = ioBundle_scan_en ? confReg_98 : confReg_82; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_99 = ioBundle_scan_en ? confReg_99 : confReg_83; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_100 = ioBundle_scan_en ? confReg_100 : confReg_84; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_101 = ioBundle_scan_en ? confReg_101 : confReg_85; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_102 = ioBundle_scan_en ? confReg_102 : confReg_86; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_103 = ioBundle_scan_en ? confReg_103 : confReg_87; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_104 = ioBundle_scan_en ? confReg_104 : confReg_88; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_105 = ioBundle_scan_en ? confReg_105 : confReg_89; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_106 = ioBundle_scan_en ? confReg_106 : confReg_90; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_107 = ioBundle_scan_en ? confReg_107 : confReg_91; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_108 = ioBundle_scan_en ? confReg_108 : confReg_92; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_109 = ioBundle_scan_en ? confReg_109 : confReg_93; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_110 = ioBundle_scan_en ? confReg_110 : confReg_94; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_111 = ioBundle_scan_en ? confReg_111 : confReg_95; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_112 = ioBundle_scan_en ? confReg_112 : confReg_96; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_113 = ioBundle_scan_en ? confReg_113 : confReg_97; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_114 = ioBundle_scan_en ? confReg_114 : confReg_98; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_115 = ioBundle_scan_en ? confReg_115 : confReg_99; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_116 = ioBundle_scan_en ? confReg_116 : confReg_100; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_117 = ioBundle_scan_en ? confReg_117 : confReg_101; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_118 = ioBundle_scan_en ? confReg_118 : confReg_102; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_119 = ioBundle_scan_en ? confReg_119 : confReg_103; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_120 = ioBundle_scan_en ? confReg_120 : confReg_104; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_121 = ioBundle_scan_en ? confReg_121 : confReg_105; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_122 = ioBundle_scan_en ? confReg_122 : confReg_106; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_123 = ioBundle_scan_en ? confReg_123 : confReg_107; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_124 = ioBundle_scan_en ? confReg_124 : confReg_108; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_125 = ioBundle_scan_en ? confReg_125 : confReg_109; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_126 = ioBundle_scan_en ? confReg_126 : confReg_110; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_127 = ioBundle_scan_en ? confReg_127 : confReg_111; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_128 = ioBundle_scan_en ? confReg_128 : confReg_112; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_129 = ioBundle_scan_en ? confReg_129 : confReg_113; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_130 = ioBundle_scan_en ? confReg_130 : confReg_114; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_131 = ioBundle_scan_en ? confReg_131 : confReg_115; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_132 = ioBundle_scan_en ? confReg_132 : confReg_116; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_133 = ioBundle_scan_en ? confReg_133 : confReg_117; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_134 = ioBundle_scan_en ? confReg_134 : confReg_118; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_135 = ioBundle_scan_en ? confReg_135 : confReg_119; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_136 = ioBundle_scan_en ? confReg_136 : confReg_120; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_137 = ioBundle_scan_en ? confReg_137 : confReg_121; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_138 = ioBundle_scan_en ? confReg_138 : confReg_122; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_139 = ioBundle_scan_en ? confReg_139 : confReg_123; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_140 = ioBundle_scan_en ? confReg_140 : confReg_124; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_141 = ioBundle_scan_en ? confReg_141 : confReg_125; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_142 = ioBundle_scan_en ? confReg_142 : confReg_126; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_143 = ioBundle_scan_en ? confReg_143 : confReg_127; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_144 = ioBundle_scan_en ? confReg_144 : confReg_128; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_145 = ioBundle_scan_en ? confReg_145 : confReg_129; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_146 = ioBundle_scan_en ? confReg_146 : confReg_130; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_147 = ioBundle_scan_en ? confReg_147 : confReg_131; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_148 = ioBundle_scan_en ? confReg_148 : confReg_132; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_149 = ioBundle_scan_en ? confReg_149 : confReg_133; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_150 = ioBundle_scan_en ? confReg_150 : confReg_134; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_151 = ioBundle_scan_en ? confReg_151 : confReg_135; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_152 = ioBundle_scan_en ? confReg_152 : confReg_136; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_153 = ioBundle_scan_en ? confReg_153 : confReg_137; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_154 = ioBundle_scan_en ? confReg_154 : confReg_138; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_155 = ioBundle_scan_en ? confReg_155 : confReg_139; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_156 = ioBundle_scan_en ? confReg_156 : confReg_140; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_157 = ioBundle_scan_en ? confReg_157 : confReg_141; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_158 = ioBundle_scan_en ? confReg_158 : confReg_142; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_159 = ioBundle_scan_en ? confReg_159 : confReg_143; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_160 = ioBundle_scan_en ? confReg_160 : confReg_144; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_161 = ioBundle_scan_en ? confReg_161 : confReg_145; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_162 = ioBundle_scan_en ? confReg_162 : confReg_146; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_163 = ioBundle_scan_en ? confReg_163 : confReg_147; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_164 = ioBundle_scan_en ? confReg_164 : confReg_148; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_165 = ioBundle_scan_en ? confReg_165 : confReg_149; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_166 = ioBundle_scan_en ? confReg_166 : confReg_150; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_167 = ioBundle_scan_en ? confReg_167 : confReg_151; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_168 = ioBundle_scan_en ? confReg_168 : confReg_152; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_169 = ioBundle_scan_en ? confReg_169 : confReg_153; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_170 = ioBundle_scan_en ? confReg_170 : confReg_154; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_171 = ioBundle_scan_en ? confReg_171 : confReg_155; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_172 = ioBundle_scan_en ? confReg_172 : confReg_156; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_173 = ioBundle_scan_en ? confReg_173 : confReg_157; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_174 = ioBundle_scan_en ? confReg_174 : confReg_158; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_175 = ioBundle_scan_en ? confReg_175 : confReg_159; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_176 = ioBundle_scan_en ? confReg_176 : confReg_160; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_177 = ioBundle_scan_en ? confReg_177 : confReg_161; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_178 = ioBundle_scan_en ? confReg_178 : confReg_162; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_179 = ioBundle_scan_en ? confReg_179 : confReg_163; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_180 = ioBundle_scan_en ? confReg_180 : confReg_164; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_181 = ioBundle_scan_en ? confReg_181 : confReg_165; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_182 = ioBundle_scan_en ? confReg_182 : confReg_166; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_183 = ioBundle_scan_en ? confReg_183 : confReg_167; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_184 = ioBundle_scan_en ? confReg_184 : confReg_168; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_185 = ioBundle_scan_en ? confReg_185 : confReg_169; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_186 = ioBundle_scan_en ? confReg_186 : confReg_170; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_187 = ioBundle_scan_en ? confReg_187 : confReg_171; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_188 = ioBundle_scan_en ? confReg_188 : confReg_172; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_189 = ioBundle_scan_en ? confReg_189 : confReg_173; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_190 = ioBundle_scan_en ? confReg_190 : confReg_174; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_191 = ioBundle_scan_en ? confReg_191 : confReg_175; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_192 = ioBundle_scan_en ? confReg_192 : confReg_176; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_193 = ioBundle_scan_en ? confReg_193 : confReg_177; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_194 = ioBundle_scan_en ? confReg_194 : confReg_178; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_195 = ioBundle_scan_en ? confReg_195 : confReg_179; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_196 = ioBundle_scan_en ? confReg_196 : confReg_180; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_197 = ioBundle_scan_en ? confReg_197 : confReg_181; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_198 = ioBundle_scan_en ? confReg_198 : confReg_182; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_199 = ioBundle_scan_en ? confReg_199 : confReg_183; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_200 = ioBundle_scan_en ? confReg_200 : confReg_184; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_201 = ioBundle_scan_en ? confReg_201 : confReg_185; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_202 = ioBundle_scan_en ? confReg_202 : confReg_186; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_203 = ioBundle_scan_en ? confReg_203 : confReg_187; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_204 = ioBundle_scan_en ? confReg_204 : confReg_188; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_205 = ioBundle_scan_en ? confReg_205 : confReg_189; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_206 = ioBundle_scan_en ? confReg_206 : confReg_190; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_207 = ioBundle_scan_en ? confReg_207 : confReg_191; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_208 = ioBundle_scan_en ? confReg_208 : confReg_192; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_209 = ioBundle_scan_en ? confReg_209 : confReg_193; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_210 = ioBundle_scan_en ? confReg_210 : confReg_194; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_211 = ioBundle_scan_en ? confReg_211 : confReg_195; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_212 = ioBundle_scan_en ? confReg_212 : confReg_196; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_213 = ioBundle_scan_en ? confReg_213 : confReg_197; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_214 = ioBundle_scan_en ? confReg_214 : confReg_198; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_215 = ioBundle_scan_en ? confReg_215 : confReg_199; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_216 = ioBundle_scan_en ? confReg_216 : confReg_200; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_217 = ioBundle_scan_en ? confReg_217 : confReg_201; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_218 = ioBundle_scan_en ? confReg_218 : confReg_202; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_219 = ioBundle_scan_en ? confReg_219 : confReg_203; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_220 = ioBundle_scan_en ? confReg_220 : confReg_204; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_221 = ioBundle_scan_en ? confReg_221 : confReg_205; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_222 = ioBundle_scan_en ? confReg_222 : confReg_206; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_223 = ioBundle_scan_en ? confReg_223 : confReg_207; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_224 = ioBundle_scan_en ? confReg_224 : confReg_208; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_225 = ioBundle_scan_en ? confReg_225 : confReg_209; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_226 = ioBundle_scan_en ? confReg_226 : confReg_210; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_227 = ioBundle_scan_en ? confReg_227 : confReg_211; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_228 = ioBundle_scan_en ? confReg_228 : confReg_212; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_229 = ioBundle_scan_en ? confReg_229 : confReg_213; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_230 = ioBundle_scan_en ? confReg_230 : confReg_214; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_231 = ioBundle_scan_en ? confReg_231 : confReg_215; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_232 = ioBundle_scan_en ? confReg_232 : confReg_216; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_233 = ioBundle_scan_en ? confReg_233 : confReg_217; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_234 = ioBundle_scan_en ? confReg_234 : confReg_218; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_235 = ioBundle_scan_en ? confReg_235 : confReg_219; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_236 = ioBundle_scan_en ? confReg_236 : confReg_220; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_237 = ioBundle_scan_en ? confReg_237 : confReg_221; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_238 = ioBundle_scan_en ? confReg_238 : confReg_222; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_239 = ioBundle_scan_en ? confReg_239 : confReg_223; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_240 = ioBundle_scan_en ? confReg_240 : confReg_224; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_241 = ioBundle_scan_en ? confReg_241 : confReg_225; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_242 = ioBundle_scan_en ? confReg_242 : confReg_226; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_243 = ioBundle_scan_en ? confReg_243 : confReg_227; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_244 = ioBundle_scan_en ? confReg_244 : confReg_228; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_245 = ioBundle_scan_en ? confReg_245 : confReg_229; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_246 = ioBundle_scan_en ? confReg_246 : confReg_230; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_247 = ioBundle_scan_en ? confReg_247 : confReg_231; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_248 = ioBundle_scan_en ? confReg_248 : confReg_232; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_249 = ioBundle_scan_en ? confReg_249 : confReg_233; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_250 = ioBundle_scan_en ? confReg_250 : confReg_234; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_251 = ioBundle_scan_en ? confReg_251 : confReg_235; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_252 = ioBundle_scan_en ? confReg_252 : confReg_236; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_253 = ioBundle_scan_en ? confReg_253 : confReg_237; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_254 = ioBundle_scan_en ? confReg_254 : confReg_238; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_255 = ioBundle_scan_en ? confReg_255 : confReg_239; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_256 = ioBundle_scan_en ? confReg_256 : confReg_240; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_257 = ioBundle_scan_en ? confReg_257 : confReg_241; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_258 = ioBundle_scan_en ? confReg_258 : confReg_242; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_259 = ioBundle_scan_en ? confReg_259 : confReg_243; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_260 = ioBundle_scan_en ? confReg_260 : confReg_244; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_261 = ioBundle_scan_en ? confReg_261 : confReg_245; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_262 = ioBundle_scan_en ? confReg_262 : confReg_246; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_263 = ioBundle_scan_en ? confReg_263 : confReg_247; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_264 = ioBundle_scan_en ? confReg_264 : confReg_248; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_265 = ioBundle_scan_en ? confReg_265 : confReg_249; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_266 = ioBundle_scan_en ? confReg_266 : confReg_250; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_267 = ioBundle_scan_en ? confReg_267 : confReg_251; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_268 = ioBundle_scan_en ? confReg_268 : confReg_252; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_269 = ioBundle_scan_en ? confReg_269 : confReg_253; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_270 = ioBundle_scan_en ? confReg_270 : confReg_254; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_271 = ioBundle_scan_en ? confReg_271 : confReg_255; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_272 = ioBundle_scan_en ? confReg_272 : confReg_256; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_273 = ioBundle_scan_en ? confReg_273 : confReg_257; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_274 = ioBundle_scan_en ? confReg_274 : confReg_258; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_275 = ioBundle_scan_en ? confReg_275 : confReg_259; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_276 = ioBundle_scan_en ? confReg_276 : confReg_260; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_277 = ioBundle_scan_en ? confReg_277 : confReg_261; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_278 = ioBundle_scan_en ? confReg_278 : confReg_262; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_279 = ioBundle_scan_en ? confReg_279 : confReg_263; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_280 = ioBundle_scan_en ? confReg_280 : confReg_264; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_281 = ioBundle_scan_en ? confReg_281 : confReg_265; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_282 = ioBundle_scan_en ? confReg_282 : confReg_266; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_283 = ioBundle_scan_en ? confReg_283 : confReg_267; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_284 = ioBundle_scan_en ? confReg_284 : confReg_268; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_285 = ioBundle_scan_en ? confReg_285 : confReg_269; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_286 = ioBundle_scan_en ? confReg_286 : confReg_270; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _GEN_287 = ioBundle_scan_en ? confReg_287 : confReg_271; // @[ScanConfRadh.scala 45:20 50:20 54:36]
  wire  _io_scan_out_WIRE_1 = confReg_1; // @[ScanConfRadh.scala 59:{25,25}]
  wire  _io_scan_out_WIRE_0 = confReg_0; // @[ScanConfRadh.scala 59:{25,25}]
  wire [1:0] io_scan_out_lo_lo_lo = {confReg_1,confReg_0}; // @[ScanConfRadh.scala 59:47]
  wire  _io_scan_out_WIRE_3 = confReg_3; // @[ScanConfRadh.scala 59:{25,25}]
  wire  _io_scan_out_WIRE_2 = confReg_2; // @[ScanConfRadh.scala 59:{25,25}]
  wire [1:0] io_scan_out_lo_lo_hi = {confReg_3,confReg_2}; // @[ScanConfRadh.scala 59:47]
  wire [3:0] io_scan_out_lo_lo = {confReg_3,confReg_2,confReg_1,confReg_0}; // @[ScanConfRadh.scala 59:47]
  wire  _io_scan_out_WIRE_5 = confReg_5; // @[ScanConfRadh.scala 59:{25,25}]
  wire  _io_scan_out_WIRE_4 = confReg_4; // @[ScanConfRadh.scala 59:{25,25}]
  wire [1:0] io_scan_out_lo_hi_lo = {confReg_5,confReg_4}; // @[ScanConfRadh.scala 59:47]
  wire  _io_scan_out_WIRE_7 = confReg_7; // @[ScanConfRadh.scala 59:{25,25}]
  wire  _io_scan_out_WIRE_6 = confReg_6; // @[ScanConfRadh.scala 59:{25,25}]
  wire [1:0] io_scan_out_lo_hi_hi = {confReg_7,confReg_6}; // @[ScanConfRadh.scala 59:47]
  wire [3:0] io_scan_out_lo_hi = {confReg_7,confReg_6,confReg_5,confReg_4}; // @[ScanConfRadh.scala 59:47]
  wire [7:0] io_scan_out_lo = {confReg_7,confReg_6,confReg_5,confReg_4,confReg_3,confReg_2,confReg_1,confReg_0}; // @[ScanConfRadh.scala 59:47]
  wire  _io_scan_out_WIRE_9 = confReg_9; // @[ScanConfRadh.scala 59:{25,25}]
  wire  _io_scan_out_WIRE_8 = confReg_8; // @[ScanConfRadh.scala 59:{25,25}]
  wire [1:0] io_scan_out_hi_lo_lo = {confReg_9,confReg_8}; // @[ScanConfRadh.scala 59:47]
  wire  _io_scan_out_WIRE_11 = confReg_11; // @[ScanConfRadh.scala 59:{25,25}]
  wire  _io_scan_out_WIRE_10 = confReg_10; // @[ScanConfRadh.scala 59:{25,25}]
  wire [1:0] io_scan_out_hi_lo_hi = {confReg_11,confReg_10}; // @[ScanConfRadh.scala 59:47]
  wire [3:0] io_scan_out_hi_lo = {confReg_11,confReg_10,confReg_9,confReg_8}; // @[ScanConfRadh.scala 59:47]
  wire  _io_scan_out_WIRE_13 = confReg_13; // @[ScanConfRadh.scala 59:{25,25}]
  wire  _io_scan_out_WIRE_12 = confReg_12; // @[ScanConfRadh.scala 59:{25,25}]
  wire [1:0] io_scan_out_hi_hi_lo = {confReg_13,confReg_12}; // @[ScanConfRadh.scala 59:47]
  wire  _io_scan_out_WIRE_15 = confReg_15; // @[ScanConfRadh.scala 59:{25,25}]
  wire  _io_scan_out_WIRE_14 = confReg_14; // @[ScanConfRadh.scala 59:{25,25}]
  wire [1:0] io_scan_out_hi_hi_hi = {confReg_15,confReg_14}; // @[ScanConfRadh.scala 59:47]
  wire [3:0] io_scan_out_hi_hi = {confReg_15,confReg_14,confReg_13,confReg_12}; // @[ScanConfRadh.scala 59:47]
  wire [7:0] io_scan_out_hi = {confReg_15,confReg_14,confReg_13,confReg_12,confReg_11,confReg_10,confReg_9,confReg_8}; // @[ScanConfRadh.scala 59:47]
  wire [15:0] io_scan_out = {confReg_15,confReg_14,confReg_13,confReg_12,confReg_11,confReg_10,confReg_9,confReg_8,
    io_scan_out_lo}; // @[ScanConfRadh.scala 59:47]
  wire  io_scan_ioLatchEnb = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 40:16 70:12]
  wire  _T = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_1 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_2 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_3 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_4 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_5 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_6 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_7 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_8 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_9 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_10 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_11 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_12 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_13 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_14 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_15 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_16 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_17 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_18 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_19 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_20 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_21 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_22 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_23 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_24 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_25 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_26 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_27 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_28 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_29 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_30 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_31 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_32 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_33 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_34 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_35 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_36 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_37 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_38 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_39 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_40 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_41 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_42 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_43 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_44 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_45 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_46 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_47 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_48 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_49 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_50 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_51 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_52 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_53 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_54 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_55 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_56 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_57 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_58 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_59 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_60 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_61 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_62 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_63 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_64 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_65 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_66 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_67 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_68 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_69 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_70 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_71 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_72 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_73 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_74 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_75 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_76 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_77 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_78 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_79 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_80 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_81 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_82 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_83 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_84 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_85 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_86 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_87 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_88 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_89 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_90 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_91 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_92 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_93 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_94 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_95 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_96 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_97 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_98 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_99 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_100 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_101 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_102 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_103 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_104 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_105 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_106 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_107 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_108 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_109 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_110 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_111 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_112 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_113 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_114 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_115 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_116 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_117 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_118 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_119 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_120 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_121 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_122 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_123 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_124 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_125 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_126 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_127 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_128 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_129 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_130 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_131 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_132 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_133 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_134 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_135 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_136 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_137 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_138 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_139 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_140 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_141 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_142 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_143 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_144 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_145 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_146 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_147 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_148 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_149 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_150 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_151 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_152 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_153 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_154 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_155 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_156 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_157 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_158 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_159 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_160 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_161 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_162 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_163 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_164 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_165 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_166 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_167 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_168 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_169 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_170 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_171 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_172 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_173 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_174 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_175 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_176 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_177 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_178 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_179 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_180 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_181 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_182 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_183 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_184 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_185 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_186 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_187 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_188 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_189 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_190 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_191 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_192 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_193 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_194 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_195 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_196 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_197 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_198 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_199 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_200 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_201 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_202 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_203 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_204 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_205 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_206 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_207 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_208 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_209 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_210 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_211 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_212 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_213 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_214 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_215 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_216 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_217 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_218 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_219 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_220 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_221 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_222 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_223 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_224 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_225 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_226 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_227 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_228 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_229 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_230 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_231 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_232 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_233 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_234 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_235 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_236 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_237 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_238 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_239 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_240 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_241 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_242 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_243 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_244 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_245 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_246 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_247 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_248 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_249 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_250 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_251 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_252 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_253 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_254 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_255 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_256 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_257 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_258 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_259 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_260 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_261 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_262 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_263 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_264 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_265 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_266 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_267 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_268 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_269 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_270 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_271 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_272 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_273 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_274 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_275 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_276 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_277 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_278 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_279 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_280 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_281 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_282 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_283 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_284 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_285 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_286 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _T_287 = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  wire  _io_confOut_WIRE_1 = b0mlcn000hn1n02x5_1_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_0 = b0mlcn000hn1n02x5_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_lo_lo_lo_lo = {_io_confOut_WIRE_1,_io_confOut_WIRE_0}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_3 = b0mlcn000hn1n02x5_3_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_2 = b0mlcn000hn1n02x5_2_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_lo_lo_lo_hi = {_io_confOut_WIRE_3,_io_confOut_WIRE_2}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_lo_lo_lo_lo_lo = {_io_confOut_WIRE_3,_io_confOut_WIRE_2,_io_confOut_WIRE_1,_io_confOut_WIRE_0
    }; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_5 = b0mlcn000hn1n02x5_5_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_4 = b0mlcn000hn1n02x5_4_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_lo_lo_hi_lo = {_io_confOut_WIRE_5,_io_confOut_WIRE_4}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_8 = b0mlcn000hn1n02x5_8_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_7 = b0mlcn000hn1n02x5_7_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_lo_lo_hi_hi_hi = {_io_confOut_WIRE_8,_io_confOut_WIRE_7}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_6 = b0mlcn000hn1n02x5_6_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_lo_lo_lo_lo_hi_hi = {_io_confOut_WIRE_8,_io_confOut_WIRE_7,_io_confOut_WIRE_6}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_lo_lo_lo_lo_hi = {_io_confOut_WIRE_8,_io_confOut_WIRE_7,_io_confOut_WIRE_6,_io_confOut_WIRE_5
    ,_io_confOut_WIRE_4}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_lo_lo_lo_lo = {_io_confOut_WIRE_8,_io_confOut_WIRE_7,_io_confOut_WIRE_6,_io_confOut_WIRE_5,
    _io_confOut_WIRE_4,_io_confOut_WIRE_3,_io_confOut_WIRE_2,_io_confOut_WIRE_1,_io_confOut_WIRE_0}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_10 = b0mlcn000hn1n02x5_10_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_9 = b0mlcn000hn1n02x5_9_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_lo_hi_lo_lo = {_io_confOut_WIRE_10,_io_confOut_WIRE_9}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_12 = b0mlcn000hn1n02x5_12_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_11 = b0mlcn000hn1n02x5_11_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_lo_hi_lo_hi = {_io_confOut_WIRE_12,_io_confOut_WIRE_11}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_lo_lo_lo_hi_lo = {_io_confOut_WIRE_12,_io_confOut_WIRE_11,_io_confOut_WIRE_10,
    _io_confOut_WIRE_9}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_14 = b0mlcn000hn1n02x5_14_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_13 = b0mlcn000hn1n02x5_13_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_lo_hi_hi_lo = {_io_confOut_WIRE_14,_io_confOut_WIRE_13}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_17 = b0mlcn000hn1n02x5_17_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_16 = b0mlcn000hn1n02x5_16_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_lo_hi_hi_hi_hi = {_io_confOut_WIRE_17,_io_confOut_WIRE_16}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_15 = b0mlcn000hn1n02x5_15_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_lo_lo_lo_hi_hi_hi = {_io_confOut_WIRE_17,_io_confOut_WIRE_16,_io_confOut_WIRE_15}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_lo_lo_lo_hi_hi = {_io_confOut_WIRE_17,_io_confOut_WIRE_16,_io_confOut_WIRE_15,
    _io_confOut_WIRE_14,_io_confOut_WIRE_13}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_lo_lo_lo_hi = {_io_confOut_WIRE_17,_io_confOut_WIRE_16,_io_confOut_WIRE_15,
    _io_confOut_WIRE_14,_io_confOut_WIRE_13,_io_confOut_WIRE_12,_io_confOut_WIRE_11,_io_confOut_WIRE_10,
    _io_confOut_WIRE_9}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_lo_lo_lo_lo = {_io_confOut_WIRE_17,_io_confOut_WIRE_16,_io_confOut_WIRE_15,_io_confOut_WIRE_14,
    _io_confOut_WIRE_13,_io_confOut_WIRE_12,_io_confOut_WIRE_11,_io_confOut_WIRE_10,_io_confOut_WIRE_9,
    io_confOut_lo_lo_lo_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_19 = b0mlcn000hn1n02x5_19_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_18 = b0mlcn000hn1n02x5_18_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_hi_lo_lo_lo = {_io_confOut_WIRE_19,_io_confOut_WIRE_18}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_21 = b0mlcn000hn1n02x5_21_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_20 = b0mlcn000hn1n02x5_20_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_hi_lo_lo_hi = {_io_confOut_WIRE_21,_io_confOut_WIRE_20}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_lo_lo_hi_lo_lo = {_io_confOut_WIRE_21,_io_confOut_WIRE_20,_io_confOut_WIRE_19,
    _io_confOut_WIRE_18}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_23 = b0mlcn000hn1n02x5_23_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_22 = b0mlcn000hn1n02x5_22_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_hi_lo_hi_lo = {_io_confOut_WIRE_23,_io_confOut_WIRE_22}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_26 = b0mlcn000hn1n02x5_26_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_25 = b0mlcn000hn1n02x5_25_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_hi_lo_hi_hi_hi = {_io_confOut_WIRE_26,_io_confOut_WIRE_25}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_24 = b0mlcn000hn1n02x5_24_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_lo_lo_hi_lo_hi_hi = {_io_confOut_WIRE_26,_io_confOut_WIRE_25,_io_confOut_WIRE_24}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_lo_lo_hi_lo_hi = {_io_confOut_WIRE_26,_io_confOut_WIRE_25,_io_confOut_WIRE_24,
    _io_confOut_WIRE_23,_io_confOut_WIRE_22}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_lo_lo_hi_lo = {_io_confOut_WIRE_26,_io_confOut_WIRE_25,_io_confOut_WIRE_24,
    _io_confOut_WIRE_23,_io_confOut_WIRE_22,_io_confOut_WIRE_21,_io_confOut_WIRE_20,_io_confOut_WIRE_19,
    _io_confOut_WIRE_18}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_28 = b0mlcn000hn1n02x5_28_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_27 = b0mlcn000hn1n02x5_27_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_hi_hi_lo_lo = {_io_confOut_WIRE_28,_io_confOut_WIRE_27}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_30 = b0mlcn000hn1n02x5_30_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_29 = b0mlcn000hn1n02x5_29_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_hi_hi_lo_hi = {_io_confOut_WIRE_30,_io_confOut_WIRE_29}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_lo_lo_hi_hi_lo = {_io_confOut_WIRE_30,_io_confOut_WIRE_29,_io_confOut_WIRE_28,
    _io_confOut_WIRE_27}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_32 = b0mlcn000hn1n02x5_32_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_31 = b0mlcn000hn1n02x5_31_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_hi_hi_hi_lo = {_io_confOut_WIRE_32,_io_confOut_WIRE_31}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_35 = b0mlcn000hn1n02x5_35_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_34 = b0mlcn000hn1n02x5_34_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_lo_hi_hi_hi_hi_hi = {_io_confOut_WIRE_35,_io_confOut_WIRE_34}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_33 = b0mlcn000hn1n02x5_33_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_lo_lo_hi_hi_hi_hi = {_io_confOut_WIRE_35,_io_confOut_WIRE_34,_io_confOut_WIRE_33}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_lo_lo_hi_hi_hi = {_io_confOut_WIRE_35,_io_confOut_WIRE_34,_io_confOut_WIRE_33,
    _io_confOut_WIRE_32,_io_confOut_WIRE_31}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_lo_lo_hi_hi = {_io_confOut_WIRE_35,_io_confOut_WIRE_34,_io_confOut_WIRE_33,
    _io_confOut_WIRE_32,_io_confOut_WIRE_31,_io_confOut_WIRE_30,_io_confOut_WIRE_29,_io_confOut_WIRE_28,
    _io_confOut_WIRE_27}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_lo_lo_lo_hi = {_io_confOut_WIRE_35,_io_confOut_WIRE_34,_io_confOut_WIRE_33,_io_confOut_WIRE_32,
    _io_confOut_WIRE_31,_io_confOut_WIRE_30,_io_confOut_WIRE_29,_io_confOut_WIRE_28,_io_confOut_WIRE_27,
    io_confOut_lo_lo_lo_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [35:0] io_confOut_lo_lo_lo = {io_confOut_lo_lo_lo_hi,io_confOut_lo_lo_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_37 = b0mlcn000hn1n02x5_37_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_36 = b0mlcn000hn1n02x5_36_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_lo_lo_lo_lo = {_io_confOut_WIRE_37,_io_confOut_WIRE_36}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_39 = b0mlcn000hn1n02x5_39_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_38 = b0mlcn000hn1n02x5_38_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_lo_lo_lo_hi = {_io_confOut_WIRE_39,_io_confOut_WIRE_38}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_lo_hi_lo_lo_lo = {_io_confOut_WIRE_39,_io_confOut_WIRE_38,_io_confOut_WIRE_37,
    _io_confOut_WIRE_36}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_41 = b0mlcn000hn1n02x5_41_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_40 = b0mlcn000hn1n02x5_40_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_lo_lo_hi_lo = {_io_confOut_WIRE_41,_io_confOut_WIRE_40}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_44 = b0mlcn000hn1n02x5_44_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_43 = b0mlcn000hn1n02x5_43_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_lo_lo_hi_hi_hi = {_io_confOut_WIRE_44,_io_confOut_WIRE_43}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_42 = b0mlcn000hn1n02x5_42_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_lo_hi_lo_lo_hi_hi = {_io_confOut_WIRE_44,_io_confOut_WIRE_43,_io_confOut_WIRE_42}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_lo_hi_lo_lo_hi = {_io_confOut_WIRE_44,_io_confOut_WIRE_43,_io_confOut_WIRE_42,
    _io_confOut_WIRE_41,_io_confOut_WIRE_40}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_lo_hi_lo_lo = {_io_confOut_WIRE_44,_io_confOut_WIRE_43,_io_confOut_WIRE_42,
    _io_confOut_WIRE_41,_io_confOut_WIRE_40,_io_confOut_WIRE_39,_io_confOut_WIRE_38,_io_confOut_WIRE_37,
    _io_confOut_WIRE_36}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_46 = b0mlcn000hn1n02x5_46_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_45 = b0mlcn000hn1n02x5_45_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_lo_hi_lo_lo = {_io_confOut_WIRE_46,_io_confOut_WIRE_45}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_48 = b0mlcn000hn1n02x5_48_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_47 = b0mlcn000hn1n02x5_47_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_lo_hi_lo_hi = {_io_confOut_WIRE_48,_io_confOut_WIRE_47}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_lo_hi_lo_hi_lo = {_io_confOut_WIRE_48,_io_confOut_WIRE_47,_io_confOut_WIRE_46,
    _io_confOut_WIRE_45}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_50 = b0mlcn000hn1n02x5_50_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_49 = b0mlcn000hn1n02x5_49_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_lo_hi_hi_lo = {_io_confOut_WIRE_50,_io_confOut_WIRE_49}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_53 = b0mlcn000hn1n02x5_53_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_52 = b0mlcn000hn1n02x5_52_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_lo_hi_hi_hi_hi = {_io_confOut_WIRE_53,_io_confOut_WIRE_52}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_51 = b0mlcn000hn1n02x5_51_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_lo_hi_lo_hi_hi_hi = {_io_confOut_WIRE_53,_io_confOut_WIRE_52,_io_confOut_WIRE_51}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_lo_hi_lo_hi_hi = {_io_confOut_WIRE_53,_io_confOut_WIRE_52,_io_confOut_WIRE_51,
    _io_confOut_WIRE_50,_io_confOut_WIRE_49}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_lo_hi_lo_hi = {_io_confOut_WIRE_53,_io_confOut_WIRE_52,_io_confOut_WIRE_51,
    _io_confOut_WIRE_50,_io_confOut_WIRE_49,_io_confOut_WIRE_48,_io_confOut_WIRE_47,_io_confOut_WIRE_46,
    _io_confOut_WIRE_45}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_lo_lo_hi_lo = {_io_confOut_WIRE_53,_io_confOut_WIRE_52,_io_confOut_WIRE_51,_io_confOut_WIRE_50,
    _io_confOut_WIRE_49,_io_confOut_WIRE_48,_io_confOut_WIRE_47,_io_confOut_WIRE_46,_io_confOut_WIRE_45,
    io_confOut_lo_lo_hi_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_55 = b0mlcn000hn1n02x5_55_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_54 = b0mlcn000hn1n02x5_54_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_hi_lo_lo_lo = {_io_confOut_WIRE_55,_io_confOut_WIRE_54}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_57 = b0mlcn000hn1n02x5_57_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_56 = b0mlcn000hn1n02x5_56_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_hi_lo_lo_hi = {_io_confOut_WIRE_57,_io_confOut_WIRE_56}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_lo_hi_hi_lo_lo = {_io_confOut_WIRE_57,_io_confOut_WIRE_56,_io_confOut_WIRE_55,
    _io_confOut_WIRE_54}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_59 = b0mlcn000hn1n02x5_59_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_58 = b0mlcn000hn1n02x5_58_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_hi_lo_hi_lo = {_io_confOut_WIRE_59,_io_confOut_WIRE_58}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_62 = b0mlcn000hn1n02x5_62_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_61 = b0mlcn000hn1n02x5_61_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_hi_lo_hi_hi_hi = {_io_confOut_WIRE_62,_io_confOut_WIRE_61}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_60 = b0mlcn000hn1n02x5_60_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_lo_hi_hi_lo_hi_hi = {_io_confOut_WIRE_62,_io_confOut_WIRE_61,_io_confOut_WIRE_60}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_lo_hi_hi_lo_hi = {_io_confOut_WIRE_62,_io_confOut_WIRE_61,_io_confOut_WIRE_60,
    _io_confOut_WIRE_59,_io_confOut_WIRE_58}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_lo_hi_hi_lo = {_io_confOut_WIRE_62,_io_confOut_WIRE_61,_io_confOut_WIRE_60,
    _io_confOut_WIRE_59,_io_confOut_WIRE_58,_io_confOut_WIRE_57,_io_confOut_WIRE_56,_io_confOut_WIRE_55,
    _io_confOut_WIRE_54}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_64 = b0mlcn000hn1n02x5_64_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_63 = b0mlcn000hn1n02x5_63_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_hi_hi_lo_lo = {_io_confOut_WIRE_64,_io_confOut_WIRE_63}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_66 = b0mlcn000hn1n02x5_66_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_65 = b0mlcn000hn1n02x5_65_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_hi_hi_lo_hi = {_io_confOut_WIRE_66,_io_confOut_WIRE_65}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_lo_hi_hi_hi_lo = {_io_confOut_WIRE_66,_io_confOut_WIRE_65,_io_confOut_WIRE_64,
    _io_confOut_WIRE_63}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_68 = b0mlcn000hn1n02x5_68_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_67 = b0mlcn000hn1n02x5_67_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_hi_hi_hi_lo = {_io_confOut_WIRE_68,_io_confOut_WIRE_67}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_71 = b0mlcn000hn1n02x5_71_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_70 = b0mlcn000hn1n02x5_70_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_lo_hi_hi_hi_hi_hi_hi = {_io_confOut_WIRE_71,_io_confOut_WIRE_70}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_69 = b0mlcn000hn1n02x5_69_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_lo_hi_hi_hi_hi_hi = {_io_confOut_WIRE_71,_io_confOut_WIRE_70,_io_confOut_WIRE_69}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_lo_hi_hi_hi_hi = {_io_confOut_WIRE_71,_io_confOut_WIRE_70,_io_confOut_WIRE_69,
    _io_confOut_WIRE_68,_io_confOut_WIRE_67}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_lo_hi_hi_hi = {_io_confOut_WIRE_71,_io_confOut_WIRE_70,_io_confOut_WIRE_69,
    _io_confOut_WIRE_68,_io_confOut_WIRE_67,_io_confOut_WIRE_66,_io_confOut_WIRE_65,_io_confOut_WIRE_64,
    _io_confOut_WIRE_63}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_lo_lo_hi_hi = {_io_confOut_WIRE_71,_io_confOut_WIRE_70,_io_confOut_WIRE_69,_io_confOut_WIRE_68,
    _io_confOut_WIRE_67,_io_confOut_WIRE_66,_io_confOut_WIRE_65,_io_confOut_WIRE_64,_io_confOut_WIRE_63,
    io_confOut_lo_lo_hi_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [35:0] io_confOut_lo_lo_hi = {io_confOut_lo_lo_hi_hi,io_confOut_lo_lo_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [71:0] io_confOut_lo_lo = {io_confOut_lo_lo_hi_hi,io_confOut_lo_lo_hi_lo,io_confOut_lo_lo_lo_hi,
    io_confOut_lo_lo_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_73 = b0mlcn000hn1n02x5_73_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_72 = b0mlcn000hn1n02x5_72_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_lo_lo_lo_lo = {_io_confOut_WIRE_73,_io_confOut_WIRE_72}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_75 = b0mlcn000hn1n02x5_75_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_74 = b0mlcn000hn1n02x5_74_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_lo_lo_lo_hi = {_io_confOut_WIRE_75,_io_confOut_WIRE_74}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_hi_lo_lo_lo_lo = {_io_confOut_WIRE_75,_io_confOut_WIRE_74,_io_confOut_WIRE_73,
    _io_confOut_WIRE_72}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_77 = b0mlcn000hn1n02x5_77_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_76 = b0mlcn000hn1n02x5_76_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_lo_lo_hi_lo = {_io_confOut_WIRE_77,_io_confOut_WIRE_76}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_80 = b0mlcn000hn1n02x5_80_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_79 = b0mlcn000hn1n02x5_79_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_lo_lo_hi_hi_hi = {_io_confOut_WIRE_80,_io_confOut_WIRE_79}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_78 = b0mlcn000hn1n02x5_78_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_hi_lo_lo_lo_hi_hi = {_io_confOut_WIRE_80,_io_confOut_WIRE_79,_io_confOut_WIRE_78}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_hi_lo_lo_lo_hi = {_io_confOut_WIRE_80,_io_confOut_WIRE_79,_io_confOut_WIRE_78,
    _io_confOut_WIRE_77,_io_confOut_WIRE_76}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_hi_lo_lo_lo = {_io_confOut_WIRE_80,_io_confOut_WIRE_79,_io_confOut_WIRE_78,
    _io_confOut_WIRE_77,_io_confOut_WIRE_76,_io_confOut_WIRE_75,_io_confOut_WIRE_74,_io_confOut_WIRE_73,
    _io_confOut_WIRE_72}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_82 = b0mlcn000hn1n02x5_82_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_81 = b0mlcn000hn1n02x5_81_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_lo_hi_lo_lo = {_io_confOut_WIRE_82,_io_confOut_WIRE_81}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_84 = b0mlcn000hn1n02x5_84_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_83 = b0mlcn000hn1n02x5_83_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_lo_hi_lo_hi = {_io_confOut_WIRE_84,_io_confOut_WIRE_83}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_hi_lo_lo_hi_lo = {_io_confOut_WIRE_84,_io_confOut_WIRE_83,_io_confOut_WIRE_82,
    _io_confOut_WIRE_81}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_86 = b0mlcn000hn1n02x5_86_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_85 = b0mlcn000hn1n02x5_85_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_lo_hi_hi_lo = {_io_confOut_WIRE_86,_io_confOut_WIRE_85}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_89 = b0mlcn000hn1n02x5_89_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_88 = b0mlcn000hn1n02x5_88_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_lo_hi_hi_hi_hi = {_io_confOut_WIRE_89,_io_confOut_WIRE_88}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_87 = b0mlcn000hn1n02x5_87_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_hi_lo_lo_hi_hi_hi = {_io_confOut_WIRE_89,_io_confOut_WIRE_88,_io_confOut_WIRE_87}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_hi_lo_lo_hi_hi = {_io_confOut_WIRE_89,_io_confOut_WIRE_88,_io_confOut_WIRE_87,
    _io_confOut_WIRE_86,_io_confOut_WIRE_85}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_hi_lo_lo_hi = {_io_confOut_WIRE_89,_io_confOut_WIRE_88,_io_confOut_WIRE_87,
    _io_confOut_WIRE_86,_io_confOut_WIRE_85,_io_confOut_WIRE_84,_io_confOut_WIRE_83,_io_confOut_WIRE_82,
    _io_confOut_WIRE_81}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_lo_hi_lo_lo = {_io_confOut_WIRE_89,_io_confOut_WIRE_88,_io_confOut_WIRE_87,_io_confOut_WIRE_86,
    _io_confOut_WIRE_85,_io_confOut_WIRE_84,_io_confOut_WIRE_83,_io_confOut_WIRE_82,_io_confOut_WIRE_81,
    io_confOut_lo_hi_lo_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_91 = b0mlcn000hn1n02x5_91_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_90 = b0mlcn000hn1n02x5_90_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_hi_lo_lo_lo = {_io_confOut_WIRE_91,_io_confOut_WIRE_90}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_93 = b0mlcn000hn1n02x5_93_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_92 = b0mlcn000hn1n02x5_92_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_hi_lo_lo_hi = {_io_confOut_WIRE_93,_io_confOut_WIRE_92}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_hi_lo_hi_lo_lo = {_io_confOut_WIRE_93,_io_confOut_WIRE_92,_io_confOut_WIRE_91,
    _io_confOut_WIRE_90}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_95 = b0mlcn000hn1n02x5_95_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_94 = b0mlcn000hn1n02x5_94_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_hi_lo_hi_lo = {_io_confOut_WIRE_95,_io_confOut_WIRE_94}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_98 = b0mlcn000hn1n02x5_98_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_97 = b0mlcn000hn1n02x5_97_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_hi_lo_hi_hi_hi = {_io_confOut_WIRE_98,_io_confOut_WIRE_97}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_96 = b0mlcn000hn1n02x5_96_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_hi_lo_hi_lo_hi_hi = {_io_confOut_WIRE_98,_io_confOut_WIRE_97,_io_confOut_WIRE_96}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_hi_lo_hi_lo_hi = {_io_confOut_WIRE_98,_io_confOut_WIRE_97,_io_confOut_WIRE_96,
    _io_confOut_WIRE_95,_io_confOut_WIRE_94}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_hi_lo_hi_lo = {_io_confOut_WIRE_98,_io_confOut_WIRE_97,_io_confOut_WIRE_96,
    _io_confOut_WIRE_95,_io_confOut_WIRE_94,_io_confOut_WIRE_93,_io_confOut_WIRE_92,_io_confOut_WIRE_91,
    _io_confOut_WIRE_90}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_100 = b0mlcn000hn1n02x5_100_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_99 = b0mlcn000hn1n02x5_99_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_hi_hi_lo_lo = {_io_confOut_WIRE_100,_io_confOut_WIRE_99}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_102 = b0mlcn000hn1n02x5_102_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_101 = b0mlcn000hn1n02x5_101_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_hi_hi_lo_hi = {_io_confOut_WIRE_102,_io_confOut_WIRE_101}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_hi_lo_hi_hi_lo = {_io_confOut_WIRE_102,_io_confOut_WIRE_101,_io_confOut_WIRE_100,
    _io_confOut_WIRE_99}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_104 = b0mlcn000hn1n02x5_104_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_103 = b0mlcn000hn1n02x5_103_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_hi_hi_hi_lo = {_io_confOut_WIRE_104,_io_confOut_WIRE_103}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_107 = b0mlcn000hn1n02x5_107_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_106 = b0mlcn000hn1n02x5_106_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_lo_hi_hi_hi_hi_hi = {_io_confOut_WIRE_107,_io_confOut_WIRE_106}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_105 = b0mlcn000hn1n02x5_105_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_hi_lo_hi_hi_hi_hi = {_io_confOut_WIRE_107,_io_confOut_WIRE_106,_io_confOut_WIRE_105}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_hi_lo_hi_hi_hi = {_io_confOut_WIRE_107,_io_confOut_WIRE_106,_io_confOut_WIRE_105,
    _io_confOut_WIRE_104,_io_confOut_WIRE_103}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_hi_lo_hi_hi = {_io_confOut_WIRE_107,_io_confOut_WIRE_106,_io_confOut_WIRE_105,
    _io_confOut_WIRE_104,_io_confOut_WIRE_103,_io_confOut_WIRE_102,_io_confOut_WIRE_101,_io_confOut_WIRE_100,
    _io_confOut_WIRE_99}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_lo_hi_lo_hi = {_io_confOut_WIRE_107,_io_confOut_WIRE_106,_io_confOut_WIRE_105,
    _io_confOut_WIRE_104,_io_confOut_WIRE_103,_io_confOut_WIRE_102,_io_confOut_WIRE_101,_io_confOut_WIRE_100,
    _io_confOut_WIRE_99,io_confOut_lo_hi_lo_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [35:0] io_confOut_lo_hi_lo = {io_confOut_lo_hi_lo_hi,io_confOut_lo_hi_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_109 = b0mlcn000hn1n02x5_109_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_108 = b0mlcn000hn1n02x5_108_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_lo_lo_lo_lo = {_io_confOut_WIRE_109,_io_confOut_WIRE_108}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_111 = b0mlcn000hn1n02x5_111_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_110 = b0mlcn000hn1n02x5_110_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_lo_lo_lo_hi = {_io_confOut_WIRE_111,_io_confOut_WIRE_110}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_hi_hi_lo_lo_lo = {_io_confOut_WIRE_111,_io_confOut_WIRE_110,_io_confOut_WIRE_109,
    _io_confOut_WIRE_108}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_113 = b0mlcn000hn1n02x5_113_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_112 = b0mlcn000hn1n02x5_112_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_lo_lo_hi_lo = {_io_confOut_WIRE_113,_io_confOut_WIRE_112}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_116 = b0mlcn000hn1n02x5_116_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_115 = b0mlcn000hn1n02x5_115_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_lo_lo_hi_hi_hi = {_io_confOut_WIRE_116,_io_confOut_WIRE_115}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_114 = b0mlcn000hn1n02x5_114_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_hi_hi_lo_lo_hi_hi = {_io_confOut_WIRE_116,_io_confOut_WIRE_115,_io_confOut_WIRE_114}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_hi_hi_lo_lo_hi = {_io_confOut_WIRE_116,_io_confOut_WIRE_115,_io_confOut_WIRE_114,
    _io_confOut_WIRE_113,_io_confOut_WIRE_112}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_hi_hi_lo_lo = {_io_confOut_WIRE_116,_io_confOut_WIRE_115,_io_confOut_WIRE_114,
    _io_confOut_WIRE_113,_io_confOut_WIRE_112,_io_confOut_WIRE_111,_io_confOut_WIRE_110,_io_confOut_WIRE_109,
    _io_confOut_WIRE_108}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_118 = b0mlcn000hn1n02x5_118_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_117 = b0mlcn000hn1n02x5_117_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_lo_hi_lo_lo = {_io_confOut_WIRE_118,_io_confOut_WIRE_117}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_120 = b0mlcn000hn1n02x5_120_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_119 = b0mlcn000hn1n02x5_119_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_lo_hi_lo_hi = {_io_confOut_WIRE_120,_io_confOut_WIRE_119}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_hi_hi_lo_hi_lo = {_io_confOut_WIRE_120,_io_confOut_WIRE_119,_io_confOut_WIRE_118,
    _io_confOut_WIRE_117}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_122 = b0mlcn000hn1n02x5_122_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_121 = b0mlcn000hn1n02x5_121_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_lo_hi_hi_lo = {_io_confOut_WIRE_122,_io_confOut_WIRE_121}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_125 = b0mlcn000hn1n02x5_125_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_124 = b0mlcn000hn1n02x5_124_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_lo_hi_hi_hi_hi = {_io_confOut_WIRE_125,_io_confOut_WIRE_124}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_123 = b0mlcn000hn1n02x5_123_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_hi_hi_lo_hi_hi_hi = {_io_confOut_WIRE_125,_io_confOut_WIRE_124,_io_confOut_WIRE_123}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_hi_hi_lo_hi_hi = {_io_confOut_WIRE_125,_io_confOut_WIRE_124,_io_confOut_WIRE_123,
    _io_confOut_WIRE_122,_io_confOut_WIRE_121}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_hi_hi_lo_hi = {_io_confOut_WIRE_125,_io_confOut_WIRE_124,_io_confOut_WIRE_123,
    _io_confOut_WIRE_122,_io_confOut_WIRE_121,_io_confOut_WIRE_120,_io_confOut_WIRE_119,_io_confOut_WIRE_118,
    _io_confOut_WIRE_117}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_lo_hi_hi_lo = {_io_confOut_WIRE_125,_io_confOut_WIRE_124,_io_confOut_WIRE_123,
    _io_confOut_WIRE_122,_io_confOut_WIRE_121,_io_confOut_WIRE_120,_io_confOut_WIRE_119,_io_confOut_WIRE_118,
    _io_confOut_WIRE_117,io_confOut_lo_hi_hi_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_127 = b0mlcn000hn1n02x5_127_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_126 = b0mlcn000hn1n02x5_126_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_hi_lo_lo_lo = {_io_confOut_WIRE_127,_io_confOut_WIRE_126}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_129 = b0mlcn000hn1n02x5_129_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_128 = b0mlcn000hn1n02x5_128_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_hi_lo_lo_hi = {_io_confOut_WIRE_129,_io_confOut_WIRE_128}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_hi_hi_hi_lo_lo = {_io_confOut_WIRE_129,_io_confOut_WIRE_128,_io_confOut_WIRE_127,
    _io_confOut_WIRE_126}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_131 = b0mlcn000hn1n02x5_131_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_130 = b0mlcn000hn1n02x5_130_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_hi_lo_hi_lo = {_io_confOut_WIRE_131,_io_confOut_WIRE_130}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_134 = b0mlcn000hn1n02x5_134_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_133 = b0mlcn000hn1n02x5_133_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_hi_lo_hi_hi_hi = {_io_confOut_WIRE_134,_io_confOut_WIRE_133}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_132 = b0mlcn000hn1n02x5_132_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_hi_hi_hi_lo_hi_hi = {_io_confOut_WIRE_134,_io_confOut_WIRE_133,_io_confOut_WIRE_132}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_hi_hi_hi_lo_hi = {_io_confOut_WIRE_134,_io_confOut_WIRE_133,_io_confOut_WIRE_132,
    _io_confOut_WIRE_131,_io_confOut_WIRE_130}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_hi_hi_hi_lo = {_io_confOut_WIRE_134,_io_confOut_WIRE_133,_io_confOut_WIRE_132,
    _io_confOut_WIRE_131,_io_confOut_WIRE_130,_io_confOut_WIRE_129,_io_confOut_WIRE_128,_io_confOut_WIRE_127,
    _io_confOut_WIRE_126}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_136 = b0mlcn000hn1n02x5_136_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_135 = b0mlcn000hn1n02x5_135_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_hi_hi_lo_lo = {_io_confOut_WIRE_136,_io_confOut_WIRE_135}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_138 = b0mlcn000hn1n02x5_138_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_137 = b0mlcn000hn1n02x5_137_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_hi_hi_lo_hi = {_io_confOut_WIRE_138,_io_confOut_WIRE_137}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_lo_hi_hi_hi_hi_lo = {_io_confOut_WIRE_138,_io_confOut_WIRE_137,_io_confOut_WIRE_136,
    _io_confOut_WIRE_135}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_140 = b0mlcn000hn1n02x5_140_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_139 = b0mlcn000hn1n02x5_139_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_hi_hi_hi_lo = {_io_confOut_WIRE_140,_io_confOut_WIRE_139}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_143 = b0mlcn000hn1n02x5_143_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_142 = b0mlcn000hn1n02x5_142_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_lo_hi_hi_hi_hi_hi_hi_hi = {_io_confOut_WIRE_143,_io_confOut_WIRE_142}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_141 = b0mlcn000hn1n02x5_141_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_lo_hi_hi_hi_hi_hi_hi = {_io_confOut_WIRE_143,_io_confOut_WIRE_142,_io_confOut_WIRE_141}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_lo_hi_hi_hi_hi_hi = {_io_confOut_WIRE_143,_io_confOut_WIRE_142,_io_confOut_WIRE_141,
    _io_confOut_WIRE_140,_io_confOut_WIRE_139}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_lo_hi_hi_hi_hi = {_io_confOut_WIRE_143,_io_confOut_WIRE_142,_io_confOut_WIRE_141,
    _io_confOut_WIRE_140,_io_confOut_WIRE_139,_io_confOut_WIRE_138,_io_confOut_WIRE_137,_io_confOut_WIRE_136,
    _io_confOut_WIRE_135}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_lo_hi_hi_hi = {_io_confOut_WIRE_143,_io_confOut_WIRE_142,_io_confOut_WIRE_141,
    _io_confOut_WIRE_140,_io_confOut_WIRE_139,_io_confOut_WIRE_138,_io_confOut_WIRE_137,_io_confOut_WIRE_136,
    _io_confOut_WIRE_135,io_confOut_lo_hi_hi_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [35:0] io_confOut_lo_hi_hi = {io_confOut_lo_hi_hi_hi,io_confOut_lo_hi_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [71:0] io_confOut_lo_hi = {io_confOut_lo_hi_hi_hi,io_confOut_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi,
    io_confOut_lo_hi_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire [143:0] io_confOut_lo = {io_confOut_lo_hi_hi_hi,io_confOut_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi,
    io_confOut_lo_hi_lo_lo,io_confOut_lo_lo_hi_hi,io_confOut_lo_lo_hi_lo,io_confOut_lo_lo_lo_hi,io_confOut_lo_lo_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_145 = b0mlcn000hn1n02x5_145_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_144 = b0mlcn000hn1n02x5_144_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_lo_lo_lo_lo = {_io_confOut_WIRE_145,_io_confOut_WIRE_144}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_147 = b0mlcn000hn1n02x5_147_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_146 = b0mlcn000hn1n02x5_146_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_lo_lo_lo_hi = {_io_confOut_WIRE_147,_io_confOut_WIRE_146}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_lo_lo_lo_lo_lo = {_io_confOut_WIRE_147,_io_confOut_WIRE_146,_io_confOut_WIRE_145,
    _io_confOut_WIRE_144}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_149 = b0mlcn000hn1n02x5_149_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_148 = b0mlcn000hn1n02x5_148_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_lo_lo_hi_lo = {_io_confOut_WIRE_149,_io_confOut_WIRE_148}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_152 = b0mlcn000hn1n02x5_152_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_151 = b0mlcn000hn1n02x5_151_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_lo_lo_hi_hi_hi = {_io_confOut_WIRE_152,_io_confOut_WIRE_151}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_150 = b0mlcn000hn1n02x5_150_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_lo_lo_lo_lo_hi_hi = {_io_confOut_WIRE_152,_io_confOut_WIRE_151,_io_confOut_WIRE_150}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_lo_lo_lo_lo_hi = {_io_confOut_WIRE_152,_io_confOut_WIRE_151,_io_confOut_WIRE_150,
    _io_confOut_WIRE_149,_io_confOut_WIRE_148}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_lo_lo_lo_lo = {_io_confOut_WIRE_152,_io_confOut_WIRE_151,_io_confOut_WIRE_150,
    _io_confOut_WIRE_149,_io_confOut_WIRE_148,_io_confOut_WIRE_147,_io_confOut_WIRE_146,_io_confOut_WIRE_145,
    _io_confOut_WIRE_144}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_154 = b0mlcn000hn1n02x5_154_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_153 = b0mlcn000hn1n02x5_153_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_lo_hi_lo_lo = {_io_confOut_WIRE_154,_io_confOut_WIRE_153}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_156 = b0mlcn000hn1n02x5_156_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_155 = b0mlcn000hn1n02x5_155_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_lo_hi_lo_hi = {_io_confOut_WIRE_156,_io_confOut_WIRE_155}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_lo_lo_lo_hi_lo = {_io_confOut_WIRE_156,_io_confOut_WIRE_155,_io_confOut_WIRE_154,
    _io_confOut_WIRE_153}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_158 = b0mlcn000hn1n02x5_158_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_157 = b0mlcn000hn1n02x5_157_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_lo_hi_hi_lo = {_io_confOut_WIRE_158,_io_confOut_WIRE_157}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_161 = b0mlcn000hn1n02x5_161_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_160 = b0mlcn000hn1n02x5_160_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_lo_hi_hi_hi_hi = {_io_confOut_WIRE_161,_io_confOut_WIRE_160}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_159 = b0mlcn000hn1n02x5_159_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_lo_lo_lo_hi_hi_hi = {_io_confOut_WIRE_161,_io_confOut_WIRE_160,_io_confOut_WIRE_159}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_lo_lo_lo_hi_hi = {_io_confOut_WIRE_161,_io_confOut_WIRE_160,_io_confOut_WIRE_159,
    _io_confOut_WIRE_158,_io_confOut_WIRE_157}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_lo_lo_lo_hi = {_io_confOut_WIRE_161,_io_confOut_WIRE_160,_io_confOut_WIRE_159,
    _io_confOut_WIRE_158,_io_confOut_WIRE_157,_io_confOut_WIRE_156,_io_confOut_WIRE_155,_io_confOut_WIRE_154,
    _io_confOut_WIRE_153}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_hi_lo_lo_lo = {_io_confOut_WIRE_161,_io_confOut_WIRE_160,_io_confOut_WIRE_159,
    _io_confOut_WIRE_158,_io_confOut_WIRE_157,_io_confOut_WIRE_156,_io_confOut_WIRE_155,_io_confOut_WIRE_154,
    _io_confOut_WIRE_153,io_confOut_hi_lo_lo_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_163 = b0mlcn000hn1n02x5_163_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_162 = b0mlcn000hn1n02x5_162_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_hi_lo_lo_lo = {_io_confOut_WIRE_163,_io_confOut_WIRE_162}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_165 = b0mlcn000hn1n02x5_165_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_164 = b0mlcn000hn1n02x5_164_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_hi_lo_lo_hi = {_io_confOut_WIRE_165,_io_confOut_WIRE_164}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_lo_lo_hi_lo_lo = {_io_confOut_WIRE_165,_io_confOut_WIRE_164,_io_confOut_WIRE_163,
    _io_confOut_WIRE_162}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_167 = b0mlcn000hn1n02x5_167_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_166 = b0mlcn000hn1n02x5_166_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_hi_lo_hi_lo = {_io_confOut_WIRE_167,_io_confOut_WIRE_166}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_170 = b0mlcn000hn1n02x5_170_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_169 = b0mlcn000hn1n02x5_169_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_hi_lo_hi_hi_hi = {_io_confOut_WIRE_170,_io_confOut_WIRE_169}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_168 = b0mlcn000hn1n02x5_168_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_lo_lo_hi_lo_hi_hi = {_io_confOut_WIRE_170,_io_confOut_WIRE_169,_io_confOut_WIRE_168}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_lo_lo_hi_lo_hi = {_io_confOut_WIRE_170,_io_confOut_WIRE_169,_io_confOut_WIRE_168,
    _io_confOut_WIRE_167,_io_confOut_WIRE_166}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_lo_lo_hi_lo = {_io_confOut_WIRE_170,_io_confOut_WIRE_169,_io_confOut_WIRE_168,
    _io_confOut_WIRE_167,_io_confOut_WIRE_166,_io_confOut_WIRE_165,_io_confOut_WIRE_164,_io_confOut_WIRE_163,
    _io_confOut_WIRE_162}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_172 = b0mlcn000hn1n02x5_172_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_171 = b0mlcn000hn1n02x5_171_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_hi_hi_lo_lo = {_io_confOut_WIRE_172,_io_confOut_WIRE_171}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_174 = b0mlcn000hn1n02x5_174_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_173 = b0mlcn000hn1n02x5_173_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_hi_hi_lo_hi = {_io_confOut_WIRE_174,_io_confOut_WIRE_173}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_lo_lo_hi_hi_lo = {_io_confOut_WIRE_174,_io_confOut_WIRE_173,_io_confOut_WIRE_172,
    _io_confOut_WIRE_171}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_176 = b0mlcn000hn1n02x5_176_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_175 = b0mlcn000hn1n02x5_175_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_hi_hi_hi_lo = {_io_confOut_WIRE_176,_io_confOut_WIRE_175}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_179 = b0mlcn000hn1n02x5_179_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_178 = b0mlcn000hn1n02x5_178_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_lo_hi_hi_hi_hi_hi = {_io_confOut_WIRE_179,_io_confOut_WIRE_178}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_177 = b0mlcn000hn1n02x5_177_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_lo_lo_hi_hi_hi_hi = {_io_confOut_WIRE_179,_io_confOut_WIRE_178,_io_confOut_WIRE_177}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_lo_lo_hi_hi_hi = {_io_confOut_WIRE_179,_io_confOut_WIRE_178,_io_confOut_WIRE_177,
    _io_confOut_WIRE_176,_io_confOut_WIRE_175}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_lo_lo_hi_hi = {_io_confOut_WIRE_179,_io_confOut_WIRE_178,_io_confOut_WIRE_177,
    _io_confOut_WIRE_176,_io_confOut_WIRE_175,_io_confOut_WIRE_174,_io_confOut_WIRE_173,_io_confOut_WIRE_172,
    _io_confOut_WIRE_171}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_hi_lo_lo_hi = {_io_confOut_WIRE_179,_io_confOut_WIRE_178,_io_confOut_WIRE_177,
    _io_confOut_WIRE_176,_io_confOut_WIRE_175,_io_confOut_WIRE_174,_io_confOut_WIRE_173,_io_confOut_WIRE_172,
    _io_confOut_WIRE_171,io_confOut_hi_lo_lo_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [35:0] io_confOut_hi_lo_lo = {io_confOut_hi_lo_lo_hi,io_confOut_hi_lo_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_181 = b0mlcn000hn1n02x5_181_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_180 = b0mlcn000hn1n02x5_180_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_lo_lo_lo_lo = {_io_confOut_WIRE_181,_io_confOut_WIRE_180}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_183 = b0mlcn000hn1n02x5_183_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_182 = b0mlcn000hn1n02x5_182_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_lo_lo_lo_hi = {_io_confOut_WIRE_183,_io_confOut_WIRE_182}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_lo_hi_lo_lo_lo = {_io_confOut_WIRE_183,_io_confOut_WIRE_182,_io_confOut_WIRE_181,
    _io_confOut_WIRE_180}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_185 = b0mlcn000hn1n02x5_185_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_184 = b0mlcn000hn1n02x5_184_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_lo_lo_hi_lo = {_io_confOut_WIRE_185,_io_confOut_WIRE_184}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_188 = b0mlcn000hn1n02x5_188_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_187 = b0mlcn000hn1n02x5_187_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_lo_lo_hi_hi_hi = {_io_confOut_WIRE_188,_io_confOut_WIRE_187}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_186 = b0mlcn000hn1n02x5_186_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_lo_hi_lo_lo_hi_hi = {_io_confOut_WIRE_188,_io_confOut_WIRE_187,_io_confOut_WIRE_186}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_lo_hi_lo_lo_hi = {_io_confOut_WIRE_188,_io_confOut_WIRE_187,_io_confOut_WIRE_186,
    _io_confOut_WIRE_185,_io_confOut_WIRE_184}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_lo_hi_lo_lo = {_io_confOut_WIRE_188,_io_confOut_WIRE_187,_io_confOut_WIRE_186,
    _io_confOut_WIRE_185,_io_confOut_WIRE_184,_io_confOut_WIRE_183,_io_confOut_WIRE_182,_io_confOut_WIRE_181,
    _io_confOut_WIRE_180}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_190 = b0mlcn000hn1n02x5_190_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_189 = b0mlcn000hn1n02x5_189_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_lo_hi_lo_lo = {_io_confOut_WIRE_190,_io_confOut_WIRE_189}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_192 = b0mlcn000hn1n02x5_192_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_191 = b0mlcn000hn1n02x5_191_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_lo_hi_lo_hi = {_io_confOut_WIRE_192,_io_confOut_WIRE_191}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_lo_hi_lo_hi_lo = {_io_confOut_WIRE_192,_io_confOut_WIRE_191,_io_confOut_WIRE_190,
    _io_confOut_WIRE_189}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_194 = b0mlcn000hn1n02x5_194_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_193 = b0mlcn000hn1n02x5_193_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_lo_hi_hi_lo = {_io_confOut_WIRE_194,_io_confOut_WIRE_193}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_197 = b0mlcn000hn1n02x5_197_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_196 = b0mlcn000hn1n02x5_196_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_lo_hi_hi_hi_hi = {_io_confOut_WIRE_197,_io_confOut_WIRE_196}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_195 = b0mlcn000hn1n02x5_195_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_lo_hi_lo_hi_hi_hi = {_io_confOut_WIRE_197,_io_confOut_WIRE_196,_io_confOut_WIRE_195}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_lo_hi_lo_hi_hi = {_io_confOut_WIRE_197,_io_confOut_WIRE_196,_io_confOut_WIRE_195,
    _io_confOut_WIRE_194,_io_confOut_WIRE_193}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_lo_hi_lo_hi = {_io_confOut_WIRE_197,_io_confOut_WIRE_196,_io_confOut_WIRE_195,
    _io_confOut_WIRE_194,_io_confOut_WIRE_193,_io_confOut_WIRE_192,_io_confOut_WIRE_191,_io_confOut_WIRE_190,
    _io_confOut_WIRE_189}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_hi_lo_hi_lo = {_io_confOut_WIRE_197,_io_confOut_WIRE_196,_io_confOut_WIRE_195,
    _io_confOut_WIRE_194,_io_confOut_WIRE_193,_io_confOut_WIRE_192,_io_confOut_WIRE_191,_io_confOut_WIRE_190,
    _io_confOut_WIRE_189,io_confOut_hi_lo_hi_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_199 = b0mlcn000hn1n02x5_199_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_198 = b0mlcn000hn1n02x5_198_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_hi_lo_lo_lo = {_io_confOut_WIRE_199,_io_confOut_WIRE_198}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_201 = b0mlcn000hn1n02x5_201_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_200 = b0mlcn000hn1n02x5_200_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_hi_lo_lo_hi = {_io_confOut_WIRE_201,_io_confOut_WIRE_200}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_lo_hi_hi_lo_lo = {_io_confOut_WIRE_201,_io_confOut_WIRE_200,_io_confOut_WIRE_199,
    _io_confOut_WIRE_198}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_203 = b0mlcn000hn1n02x5_203_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_202 = b0mlcn000hn1n02x5_202_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_hi_lo_hi_lo = {_io_confOut_WIRE_203,_io_confOut_WIRE_202}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_206 = b0mlcn000hn1n02x5_206_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_205 = b0mlcn000hn1n02x5_205_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_hi_lo_hi_hi_hi = {_io_confOut_WIRE_206,_io_confOut_WIRE_205}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_204 = b0mlcn000hn1n02x5_204_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_lo_hi_hi_lo_hi_hi = {_io_confOut_WIRE_206,_io_confOut_WIRE_205,_io_confOut_WIRE_204}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_lo_hi_hi_lo_hi = {_io_confOut_WIRE_206,_io_confOut_WIRE_205,_io_confOut_WIRE_204,
    _io_confOut_WIRE_203,_io_confOut_WIRE_202}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_lo_hi_hi_lo = {_io_confOut_WIRE_206,_io_confOut_WIRE_205,_io_confOut_WIRE_204,
    _io_confOut_WIRE_203,_io_confOut_WIRE_202,_io_confOut_WIRE_201,_io_confOut_WIRE_200,_io_confOut_WIRE_199,
    _io_confOut_WIRE_198}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_208 = b0mlcn000hn1n02x5_208_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_207 = b0mlcn000hn1n02x5_207_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_hi_hi_lo_lo = {_io_confOut_WIRE_208,_io_confOut_WIRE_207}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_210 = b0mlcn000hn1n02x5_210_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_209 = b0mlcn000hn1n02x5_209_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_hi_hi_lo_hi = {_io_confOut_WIRE_210,_io_confOut_WIRE_209}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_lo_hi_hi_hi_lo = {_io_confOut_WIRE_210,_io_confOut_WIRE_209,_io_confOut_WIRE_208,
    _io_confOut_WIRE_207}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_212 = b0mlcn000hn1n02x5_212_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_211 = b0mlcn000hn1n02x5_211_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_hi_hi_hi_lo = {_io_confOut_WIRE_212,_io_confOut_WIRE_211}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_215 = b0mlcn000hn1n02x5_215_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_214 = b0mlcn000hn1n02x5_214_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_lo_hi_hi_hi_hi_hi_hi = {_io_confOut_WIRE_215,_io_confOut_WIRE_214}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_213 = b0mlcn000hn1n02x5_213_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_lo_hi_hi_hi_hi_hi = {_io_confOut_WIRE_215,_io_confOut_WIRE_214,_io_confOut_WIRE_213}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_lo_hi_hi_hi_hi = {_io_confOut_WIRE_215,_io_confOut_WIRE_214,_io_confOut_WIRE_213,
    _io_confOut_WIRE_212,_io_confOut_WIRE_211}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_lo_hi_hi_hi = {_io_confOut_WIRE_215,_io_confOut_WIRE_214,_io_confOut_WIRE_213,
    _io_confOut_WIRE_212,_io_confOut_WIRE_211,_io_confOut_WIRE_210,_io_confOut_WIRE_209,_io_confOut_WIRE_208,
    _io_confOut_WIRE_207}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_hi_lo_hi_hi = {_io_confOut_WIRE_215,_io_confOut_WIRE_214,_io_confOut_WIRE_213,
    _io_confOut_WIRE_212,_io_confOut_WIRE_211,_io_confOut_WIRE_210,_io_confOut_WIRE_209,_io_confOut_WIRE_208,
    _io_confOut_WIRE_207,io_confOut_hi_lo_hi_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [35:0] io_confOut_hi_lo_hi = {io_confOut_hi_lo_hi_hi,io_confOut_hi_lo_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [71:0] io_confOut_hi_lo = {io_confOut_hi_lo_hi_hi,io_confOut_hi_lo_hi_lo,io_confOut_hi_lo_lo_hi,
    io_confOut_hi_lo_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_217 = b0mlcn000hn1n02x5_217_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_216 = b0mlcn000hn1n02x5_216_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_lo_lo_lo_lo = {_io_confOut_WIRE_217,_io_confOut_WIRE_216}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_219 = b0mlcn000hn1n02x5_219_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_218 = b0mlcn000hn1n02x5_218_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_lo_lo_lo_hi = {_io_confOut_WIRE_219,_io_confOut_WIRE_218}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_hi_lo_lo_lo_lo = {_io_confOut_WIRE_219,_io_confOut_WIRE_218,_io_confOut_WIRE_217,
    _io_confOut_WIRE_216}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_221 = b0mlcn000hn1n02x5_221_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_220 = b0mlcn000hn1n02x5_220_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_lo_lo_hi_lo = {_io_confOut_WIRE_221,_io_confOut_WIRE_220}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_224 = b0mlcn000hn1n02x5_224_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_223 = b0mlcn000hn1n02x5_223_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_lo_lo_hi_hi_hi = {_io_confOut_WIRE_224,_io_confOut_WIRE_223}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_222 = b0mlcn000hn1n02x5_222_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_hi_lo_lo_lo_hi_hi = {_io_confOut_WIRE_224,_io_confOut_WIRE_223,_io_confOut_WIRE_222}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_hi_lo_lo_lo_hi = {_io_confOut_WIRE_224,_io_confOut_WIRE_223,_io_confOut_WIRE_222,
    _io_confOut_WIRE_221,_io_confOut_WIRE_220}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_hi_lo_lo_lo = {_io_confOut_WIRE_224,_io_confOut_WIRE_223,_io_confOut_WIRE_222,
    _io_confOut_WIRE_221,_io_confOut_WIRE_220,_io_confOut_WIRE_219,_io_confOut_WIRE_218,_io_confOut_WIRE_217,
    _io_confOut_WIRE_216}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_226 = b0mlcn000hn1n02x5_226_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_225 = b0mlcn000hn1n02x5_225_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_lo_hi_lo_lo = {_io_confOut_WIRE_226,_io_confOut_WIRE_225}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_228 = b0mlcn000hn1n02x5_228_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_227 = b0mlcn000hn1n02x5_227_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_lo_hi_lo_hi = {_io_confOut_WIRE_228,_io_confOut_WIRE_227}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_hi_lo_lo_hi_lo = {_io_confOut_WIRE_228,_io_confOut_WIRE_227,_io_confOut_WIRE_226,
    _io_confOut_WIRE_225}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_230 = b0mlcn000hn1n02x5_230_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_229 = b0mlcn000hn1n02x5_229_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_lo_hi_hi_lo = {_io_confOut_WIRE_230,_io_confOut_WIRE_229}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_233 = b0mlcn000hn1n02x5_233_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_232 = b0mlcn000hn1n02x5_232_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_lo_hi_hi_hi_hi = {_io_confOut_WIRE_233,_io_confOut_WIRE_232}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_231 = b0mlcn000hn1n02x5_231_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_hi_lo_lo_hi_hi_hi = {_io_confOut_WIRE_233,_io_confOut_WIRE_232,_io_confOut_WIRE_231}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_hi_lo_lo_hi_hi = {_io_confOut_WIRE_233,_io_confOut_WIRE_232,_io_confOut_WIRE_231,
    _io_confOut_WIRE_230,_io_confOut_WIRE_229}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_hi_lo_lo_hi = {_io_confOut_WIRE_233,_io_confOut_WIRE_232,_io_confOut_WIRE_231,
    _io_confOut_WIRE_230,_io_confOut_WIRE_229,_io_confOut_WIRE_228,_io_confOut_WIRE_227,_io_confOut_WIRE_226,
    _io_confOut_WIRE_225}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_hi_hi_lo_lo = {_io_confOut_WIRE_233,_io_confOut_WIRE_232,_io_confOut_WIRE_231,
    _io_confOut_WIRE_230,_io_confOut_WIRE_229,_io_confOut_WIRE_228,_io_confOut_WIRE_227,_io_confOut_WIRE_226,
    _io_confOut_WIRE_225,io_confOut_hi_hi_lo_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_235 = b0mlcn000hn1n02x5_235_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_234 = b0mlcn000hn1n02x5_234_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_hi_lo_lo_lo = {_io_confOut_WIRE_235,_io_confOut_WIRE_234}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_237 = b0mlcn000hn1n02x5_237_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_236 = b0mlcn000hn1n02x5_236_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_hi_lo_lo_hi = {_io_confOut_WIRE_237,_io_confOut_WIRE_236}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_hi_lo_hi_lo_lo = {_io_confOut_WIRE_237,_io_confOut_WIRE_236,_io_confOut_WIRE_235,
    _io_confOut_WIRE_234}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_239 = b0mlcn000hn1n02x5_239_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_238 = b0mlcn000hn1n02x5_238_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_hi_lo_hi_lo = {_io_confOut_WIRE_239,_io_confOut_WIRE_238}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_242 = b0mlcn000hn1n02x5_242_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_241 = b0mlcn000hn1n02x5_241_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_hi_lo_hi_hi_hi = {_io_confOut_WIRE_242,_io_confOut_WIRE_241}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_240 = b0mlcn000hn1n02x5_240_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_hi_lo_hi_lo_hi_hi = {_io_confOut_WIRE_242,_io_confOut_WIRE_241,_io_confOut_WIRE_240}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_hi_lo_hi_lo_hi = {_io_confOut_WIRE_242,_io_confOut_WIRE_241,_io_confOut_WIRE_240,
    _io_confOut_WIRE_239,_io_confOut_WIRE_238}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_hi_lo_hi_lo = {_io_confOut_WIRE_242,_io_confOut_WIRE_241,_io_confOut_WIRE_240,
    _io_confOut_WIRE_239,_io_confOut_WIRE_238,_io_confOut_WIRE_237,_io_confOut_WIRE_236,_io_confOut_WIRE_235,
    _io_confOut_WIRE_234}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_244 = b0mlcn000hn1n02x5_244_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_243 = b0mlcn000hn1n02x5_243_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_hi_hi_lo_lo = {_io_confOut_WIRE_244,_io_confOut_WIRE_243}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_246 = b0mlcn000hn1n02x5_246_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_245 = b0mlcn000hn1n02x5_245_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_hi_hi_lo_hi = {_io_confOut_WIRE_246,_io_confOut_WIRE_245}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_hi_lo_hi_hi_lo = {_io_confOut_WIRE_246,_io_confOut_WIRE_245,_io_confOut_WIRE_244,
    _io_confOut_WIRE_243}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_248 = b0mlcn000hn1n02x5_248_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_247 = b0mlcn000hn1n02x5_247_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_hi_hi_hi_lo = {_io_confOut_WIRE_248,_io_confOut_WIRE_247}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_251 = b0mlcn000hn1n02x5_251_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_250 = b0mlcn000hn1n02x5_250_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_lo_hi_hi_hi_hi_hi = {_io_confOut_WIRE_251,_io_confOut_WIRE_250}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_249 = b0mlcn000hn1n02x5_249_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_hi_lo_hi_hi_hi_hi = {_io_confOut_WIRE_251,_io_confOut_WIRE_250,_io_confOut_WIRE_249}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_hi_lo_hi_hi_hi = {_io_confOut_WIRE_251,_io_confOut_WIRE_250,_io_confOut_WIRE_249,
    _io_confOut_WIRE_248,_io_confOut_WIRE_247}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_hi_lo_hi_hi = {_io_confOut_WIRE_251,_io_confOut_WIRE_250,_io_confOut_WIRE_249,
    _io_confOut_WIRE_248,_io_confOut_WIRE_247,_io_confOut_WIRE_246,_io_confOut_WIRE_245,_io_confOut_WIRE_244,
    _io_confOut_WIRE_243}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_hi_hi_lo_hi = {_io_confOut_WIRE_251,_io_confOut_WIRE_250,_io_confOut_WIRE_249,
    _io_confOut_WIRE_248,_io_confOut_WIRE_247,_io_confOut_WIRE_246,_io_confOut_WIRE_245,_io_confOut_WIRE_244,
    _io_confOut_WIRE_243,io_confOut_hi_hi_lo_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [35:0] io_confOut_hi_hi_lo = {io_confOut_hi_hi_lo_hi,io_confOut_hi_hi_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_253 = b0mlcn000hn1n02x5_253_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_252 = b0mlcn000hn1n02x5_252_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_lo_lo_lo_lo = {_io_confOut_WIRE_253,_io_confOut_WIRE_252}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_255 = b0mlcn000hn1n02x5_255_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_254 = b0mlcn000hn1n02x5_254_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_lo_lo_lo_hi = {_io_confOut_WIRE_255,_io_confOut_WIRE_254}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_hi_hi_lo_lo_lo = {_io_confOut_WIRE_255,_io_confOut_WIRE_254,_io_confOut_WIRE_253,
    _io_confOut_WIRE_252}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_257 = b0mlcn000hn1n02x5_257_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_256 = b0mlcn000hn1n02x5_256_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_lo_lo_hi_lo = {_io_confOut_WIRE_257,_io_confOut_WIRE_256}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_260 = b0mlcn000hn1n02x5_260_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_259 = b0mlcn000hn1n02x5_259_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_lo_lo_hi_hi_hi = {_io_confOut_WIRE_260,_io_confOut_WIRE_259}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_258 = b0mlcn000hn1n02x5_258_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_hi_hi_lo_lo_hi_hi = {_io_confOut_WIRE_260,_io_confOut_WIRE_259,_io_confOut_WIRE_258}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_hi_hi_lo_lo_hi = {_io_confOut_WIRE_260,_io_confOut_WIRE_259,_io_confOut_WIRE_258,
    _io_confOut_WIRE_257,_io_confOut_WIRE_256}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_hi_hi_lo_lo = {_io_confOut_WIRE_260,_io_confOut_WIRE_259,_io_confOut_WIRE_258,
    _io_confOut_WIRE_257,_io_confOut_WIRE_256,_io_confOut_WIRE_255,_io_confOut_WIRE_254,_io_confOut_WIRE_253,
    _io_confOut_WIRE_252}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_262 = b0mlcn000hn1n02x5_262_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_261 = b0mlcn000hn1n02x5_261_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_lo_hi_lo_lo = {_io_confOut_WIRE_262,_io_confOut_WIRE_261}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_264 = b0mlcn000hn1n02x5_264_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_263 = b0mlcn000hn1n02x5_263_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_lo_hi_lo_hi = {_io_confOut_WIRE_264,_io_confOut_WIRE_263}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_hi_hi_lo_hi_lo = {_io_confOut_WIRE_264,_io_confOut_WIRE_263,_io_confOut_WIRE_262,
    _io_confOut_WIRE_261}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_266 = b0mlcn000hn1n02x5_266_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_265 = b0mlcn000hn1n02x5_265_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_lo_hi_hi_lo = {_io_confOut_WIRE_266,_io_confOut_WIRE_265}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_269 = b0mlcn000hn1n02x5_269_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_268 = b0mlcn000hn1n02x5_268_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_lo_hi_hi_hi_hi = {_io_confOut_WIRE_269,_io_confOut_WIRE_268}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_267 = b0mlcn000hn1n02x5_267_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_hi_hi_lo_hi_hi_hi = {_io_confOut_WIRE_269,_io_confOut_WIRE_268,_io_confOut_WIRE_267}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_hi_hi_lo_hi_hi = {_io_confOut_WIRE_269,_io_confOut_WIRE_268,_io_confOut_WIRE_267,
    _io_confOut_WIRE_266,_io_confOut_WIRE_265}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_hi_hi_lo_hi = {_io_confOut_WIRE_269,_io_confOut_WIRE_268,_io_confOut_WIRE_267,
    _io_confOut_WIRE_266,_io_confOut_WIRE_265,_io_confOut_WIRE_264,_io_confOut_WIRE_263,_io_confOut_WIRE_262,
    _io_confOut_WIRE_261}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_hi_hi_hi_lo = {_io_confOut_WIRE_269,_io_confOut_WIRE_268,_io_confOut_WIRE_267,
    _io_confOut_WIRE_266,_io_confOut_WIRE_265,_io_confOut_WIRE_264,_io_confOut_WIRE_263,_io_confOut_WIRE_262,
    _io_confOut_WIRE_261,io_confOut_hi_hi_hi_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_271 = b0mlcn000hn1n02x5_271_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_270 = b0mlcn000hn1n02x5_270_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_hi_lo_lo_lo = {_io_confOut_WIRE_271,_io_confOut_WIRE_270}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_273 = b0mlcn000hn1n02x5_273_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_272 = b0mlcn000hn1n02x5_272_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_hi_lo_lo_hi = {_io_confOut_WIRE_273,_io_confOut_WIRE_272}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_hi_hi_hi_lo_lo = {_io_confOut_WIRE_273,_io_confOut_WIRE_272,_io_confOut_WIRE_271,
    _io_confOut_WIRE_270}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_275 = b0mlcn000hn1n02x5_275_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_274 = b0mlcn000hn1n02x5_274_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_hi_lo_hi_lo = {_io_confOut_WIRE_275,_io_confOut_WIRE_274}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_278 = b0mlcn000hn1n02x5_278_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_277 = b0mlcn000hn1n02x5_277_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_hi_lo_hi_hi_hi = {_io_confOut_WIRE_278,_io_confOut_WIRE_277}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_276 = b0mlcn000hn1n02x5_276_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_hi_hi_hi_lo_hi_hi = {_io_confOut_WIRE_278,_io_confOut_WIRE_277,_io_confOut_WIRE_276}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_hi_hi_hi_lo_hi = {_io_confOut_WIRE_278,_io_confOut_WIRE_277,_io_confOut_WIRE_276,
    _io_confOut_WIRE_275,_io_confOut_WIRE_274}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_hi_hi_hi_lo = {_io_confOut_WIRE_278,_io_confOut_WIRE_277,_io_confOut_WIRE_276,
    _io_confOut_WIRE_275,_io_confOut_WIRE_274,_io_confOut_WIRE_273,_io_confOut_WIRE_272,_io_confOut_WIRE_271,
    _io_confOut_WIRE_270}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_280 = b0mlcn000hn1n02x5_280_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_279 = b0mlcn000hn1n02x5_279_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_hi_hi_lo_lo = {_io_confOut_WIRE_280,_io_confOut_WIRE_279}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_282 = b0mlcn000hn1n02x5_282_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_281 = b0mlcn000hn1n02x5_281_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_hi_hi_lo_hi = {_io_confOut_WIRE_282,_io_confOut_WIRE_281}; // @[ScanConfRadh.scala 67:45]
  wire [3:0] io_confOut_hi_hi_hi_hi_hi_lo = {_io_confOut_WIRE_282,_io_confOut_WIRE_281,_io_confOut_WIRE_280,
    _io_confOut_WIRE_279}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_284 = b0mlcn000hn1n02x5_284_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_283 = b0mlcn000hn1n02x5_283_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_hi_hi_hi_lo = {_io_confOut_WIRE_284,_io_confOut_WIRE_283}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_287 = b0mlcn000hn1n02x5_287_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire  _io_confOut_WIRE_286 = b0mlcn000hn1n02x5_286_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [1:0] io_confOut_hi_hi_hi_hi_hi_hi_hi_hi = {_io_confOut_WIRE_287,_io_confOut_WIRE_286}; // @[ScanConfRadh.scala 67:45]
  wire  _io_confOut_WIRE_285 = b0mlcn000hn1n02x5_285_o; // @[ScanConfRadh.scala 67:{24,24}]
  wire [2:0] io_confOut_hi_hi_hi_hi_hi_hi_hi = {_io_confOut_WIRE_287,_io_confOut_WIRE_286,_io_confOut_WIRE_285}; // @[ScanConfRadh.scala 67:45]
  wire [4:0] io_confOut_hi_hi_hi_hi_hi_hi = {_io_confOut_WIRE_287,_io_confOut_WIRE_286,_io_confOut_WIRE_285,
    _io_confOut_WIRE_284,_io_confOut_WIRE_283}; // @[ScanConfRadh.scala 67:45]
  wire [8:0] io_confOut_hi_hi_hi_hi_hi = {_io_confOut_WIRE_287,_io_confOut_WIRE_286,_io_confOut_WIRE_285,
    _io_confOut_WIRE_284,_io_confOut_WIRE_283,_io_confOut_WIRE_282,_io_confOut_WIRE_281,_io_confOut_WIRE_280,
    _io_confOut_WIRE_279}; // @[ScanConfRadh.scala 67:45]
  wire [17:0] io_confOut_hi_hi_hi_hi = {_io_confOut_WIRE_287,_io_confOut_WIRE_286,_io_confOut_WIRE_285,
    _io_confOut_WIRE_284,_io_confOut_WIRE_283,_io_confOut_WIRE_282,_io_confOut_WIRE_281,_io_confOut_WIRE_280,
    _io_confOut_WIRE_279,io_confOut_hi_hi_hi_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [35:0] io_confOut_hi_hi_hi = {io_confOut_hi_hi_hi_hi,io_confOut_hi_hi_hi_lo}; // @[ScanConfRadh.scala 67:45]
  wire [71:0] io_confOut_hi_hi = {io_confOut_hi_hi_hi_hi,io_confOut_hi_hi_hi_lo,io_confOut_hi_hi_lo_hi,
    io_confOut_hi_hi_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire [143:0] io_confOut_hi = {io_confOut_hi_hi_hi_hi,io_confOut_hi_hi_hi_lo,io_confOut_hi_hi_lo_hi,
    io_confOut_hi_hi_lo_lo,io_confOut_hi_lo_hi_hi,io_confOut_hi_lo_hi_lo,io_confOut_hi_lo_lo_hi,io_confOut_hi_lo_lo_lo}; // @[ScanConfRadh.scala 67:45]
  wire [287:0] io_confOut = {io_confOut_hi_hi_hi_hi,io_confOut_hi_hi_hi_lo,io_confOut_hi_hi_lo_hi,io_confOut_hi_hi_lo_lo
    ,io_confOut_hi_lo_hi_hi,io_confOut_hi_lo_hi_lo,io_confOut_hi_lo_lo_hi,io_confOut_hi_lo_lo_lo,io_confOut_lo}; // @[ScanConfRadh.scala 67:45]
  wire [287:0] _io_confOut_T = io_confOut; // @[ScanConfRadh.scala 67:45]
  wire [15:0] _io_scan_out_T = io_scan_out; // @[ScanConfRadh.scala 59:47]
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_d),
    .clk(b0mlcn000hn1n02x5_clk),
    .o(b0mlcn000hn1n02x5_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_1 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_1_d),
    .clk(b0mlcn000hn1n02x5_1_clk),
    .o(b0mlcn000hn1n02x5_1_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_2 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_2_d),
    .clk(b0mlcn000hn1n02x5_2_clk),
    .o(b0mlcn000hn1n02x5_2_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_3 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_3_d),
    .clk(b0mlcn000hn1n02x5_3_clk),
    .o(b0mlcn000hn1n02x5_3_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_4 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_4_d),
    .clk(b0mlcn000hn1n02x5_4_clk),
    .o(b0mlcn000hn1n02x5_4_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_5 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_5_d),
    .clk(b0mlcn000hn1n02x5_5_clk),
    .o(b0mlcn000hn1n02x5_5_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_6 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_6_d),
    .clk(b0mlcn000hn1n02x5_6_clk),
    .o(b0mlcn000hn1n02x5_6_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_7 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_7_d),
    .clk(b0mlcn000hn1n02x5_7_clk),
    .o(b0mlcn000hn1n02x5_7_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_8 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_8_d),
    .clk(b0mlcn000hn1n02x5_8_clk),
    .o(b0mlcn000hn1n02x5_8_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_9 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_9_d),
    .clk(b0mlcn000hn1n02x5_9_clk),
    .o(b0mlcn000hn1n02x5_9_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_10 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_10_d),
    .clk(b0mlcn000hn1n02x5_10_clk),
    .o(b0mlcn000hn1n02x5_10_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_11 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_11_d),
    .clk(b0mlcn000hn1n02x5_11_clk),
    .o(b0mlcn000hn1n02x5_11_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_12 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_12_d),
    .clk(b0mlcn000hn1n02x5_12_clk),
    .o(b0mlcn000hn1n02x5_12_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_13 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_13_d),
    .clk(b0mlcn000hn1n02x5_13_clk),
    .o(b0mlcn000hn1n02x5_13_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_14 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_14_d),
    .clk(b0mlcn000hn1n02x5_14_clk),
    .o(b0mlcn000hn1n02x5_14_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_15 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_15_d),
    .clk(b0mlcn000hn1n02x5_15_clk),
    .o(b0mlcn000hn1n02x5_15_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_16 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_16_d),
    .clk(b0mlcn000hn1n02x5_16_clk),
    .o(b0mlcn000hn1n02x5_16_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_17 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_17_d),
    .clk(b0mlcn000hn1n02x5_17_clk),
    .o(b0mlcn000hn1n02x5_17_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_18 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_18_d),
    .clk(b0mlcn000hn1n02x5_18_clk),
    .o(b0mlcn000hn1n02x5_18_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_19 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_19_d),
    .clk(b0mlcn000hn1n02x5_19_clk),
    .o(b0mlcn000hn1n02x5_19_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_20 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_20_d),
    .clk(b0mlcn000hn1n02x5_20_clk),
    .o(b0mlcn000hn1n02x5_20_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_21 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_21_d),
    .clk(b0mlcn000hn1n02x5_21_clk),
    .o(b0mlcn000hn1n02x5_21_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_22 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_22_d),
    .clk(b0mlcn000hn1n02x5_22_clk),
    .o(b0mlcn000hn1n02x5_22_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_23 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_23_d),
    .clk(b0mlcn000hn1n02x5_23_clk),
    .o(b0mlcn000hn1n02x5_23_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_24 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_24_d),
    .clk(b0mlcn000hn1n02x5_24_clk),
    .o(b0mlcn000hn1n02x5_24_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_25 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_25_d),
    .clk(b0mlcn000hn1n02x5_25_clk),
    .o(b0mlcn000hn1n02x5_25_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_26 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_26_d),
    .clk(b0mlcn000hn1n02x5_26_clk),
    .o(b0mlcn000hn1n02x5_26_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_27 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_27_d),
    .clk(b0mlcn000hn1n02x5_27_clk),
    .o(b0mlcn000hn1n02x5_27_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_28 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_28_d),
    .clk(b0mlcn000hn1n02x5_28_clk),
    .o(b0mlcn000hn1n02x5_28_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_29 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_29_d),
    .clk(b0mlcn000hn1n02x5_29_clk),
    .o(b0mlcn000hn1n02x5_29_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_30 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_30_d),
    .clk(b0mlcn000hn1n02x5_30_clk),
    .o(b0mlcn000hn1n02x5_30_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_31 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_31_d),
    .clk(b0mlcn000hn1n02x5_31_clk),
    .o(b0mlcn000hn1n02x5_31_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_32 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_32_d),
    .clk(b0mlcn000hn1n02x5_32_clk),
    .o(b0mlcn000hn1n02x5_32_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_33 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_33_d),
    .clk(b0mlcn000hn1n02x5_33_clk),
    .o(b0mlcn000hn1n02x5_33_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_34 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_34_d),
    .clk(b0mlcn000hn1n02x5_34_clk),
    .o(b0mlcn000hn1n02x5_34_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_35 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_35_d),
    .clk(b0mlcn000hn1n02x5_35_clk),
    .o(b0mlcn000hn1n02x5_35_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_36 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_36_d),
    .clk(b0mlcn000hn1n02x5_36_clk),
    .o(b0mlcn000hn1n02x5_36_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_37 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_37_d),
    .clk(b0mlcn000hn1n02x5_37_clk),
    .o(b0mlcn000hn1n02x5_37_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_38 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_38_d),
    .clk(b0mlcn000hn1n02x5_38_clk),
    .o(b0mlcn000hn1n02x5_38_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_39 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_39_d),
    .clk(b0mlcn000hn1n02x5_39_clk),
    .o(b0mlcn000hn1n02x5_39_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_40 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_40_d),
    .clk(b0mlcn000hn1n02x5_40_clk),
    .o(b0mlcn000hn1n02x5_40_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_41 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_41_d),
    .clk(b0mlcn000hn1n02x5_41_clk),
    .o(b0mlcn000hn1n02x5_41_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_42 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_42_d),
    .clk(b0mlcn000hn1n02x5_42_clk),
    .o(b0mlcn000hn1n02x5_42_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_43 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_43_d),
    .clk(b0mlcn000hn1n02x5_43_clk),
    .o(b0mlcn000hn1n02x5_43_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_44 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_44_d),
    .clk(b0mlcn000hn1n02x5_44_clk),
    .o(b0mlcn000hn1n02x5_44_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_45 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_45_d),
    .clk(b0mlcn000hn1n02x5_45_clk),
    .o(b0mlcn000hn1n02x5_45_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_46 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_46_d),
    .clk(b0mlcn000hn1n02x5_46_clk),
    .o(b0mlcn000hn1n02x5_46_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_47 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_47_d),
    .clk(b0mlcn000hn1n02x5_47_clk),
    .o(b0mlcn000hn1n02x5_47_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_48 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_48_d),
    .clk(b0mlcn000hn1n02x5_48_clk),
    .o(b0mlcn000hn1n02x5_48_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_49 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_49_d),
    .clk(b0mlcn000hn1n02x5_49_clk),
    .o(b0mlcn000hn1n02x5_49_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_50 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_50_d),
    .clk(b0mlcn000hn1n02x5_50_clk),
    .o(b0mlcn000hn1n02x5_50_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_51 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_51_d),
    .clk(b0mlcn000hn1n02x5_51_clk),
    .o(b0mlcn000hn1n02x5_51_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_52 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_52_d),
    .clk(b0mlcn000hn1n02x5_52_clk),
    .o(b0mlcn000hn1n02x5_52_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_53 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_53_d),
    .clk(b0mlcn000hn1n02x5_53_clk),
    .o(b0mlcn000hn1n02x5_53_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_54 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_54_d),
    .clk(b0mlcn000hn1n02x5_54_clk),
    .o(b0mlcn000hn1n02x5_54_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_55 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_55_d),
    .clk(b0mlcn000hn1n02x5_55_clk),
    .o(b0mlcn000hn1n02x5_55_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_56 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_56_d),
    .clk(b0mlcn000hn1n02x5_56_clk),
    .o(b0mlcn000hn1n02x5_56_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_57 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_57_d),
    .clk(b0mlcn000hn1n02x5_57_clk),
    .o(b0mlcn000hn1n02x5_57_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_58 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_58_d),
    .clk(b0mlcn000hn1n02x5_58_clk),
    .o(b0mlcn000hn1n02x5_58_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_59 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_59_d),
    .clk(b0mlcn000hn1n02x5_59_clk),
    .o(b0mlcn000hn1n02x5_59_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_60 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_60_d),
    .clk(b0mlcn000hn1n02x5_60_clk),
    .o(b0mlcn000hn1n02x5_60_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_61 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_61_d),
    .clk(b0mlcn000hn1n02x5_61_clk),
    .o(b0mlcn000hn1n02x5_61_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_62 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_62_d),
    .clk(b0mlcn000hn1n02x5_62_clk),
    .o(b0mlcn000hn1n02x5_62_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_63 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_63_d),
    .clk(b0mlcn000hn1n02x5_63_clk),
    .o(b0mlcn000hn1n02x5_63_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_64 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_64_d),
    .clk(b0mlcn000hn1n02x5_64_clk),
    .o(b0mlcn000hn1n02x5_64_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_65 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_65_d),
    .clk(b0mlcn000hn1n02x5_65_clk),
    .o(b0mlcn000hn1n02x5_65_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_66 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_66_d),
    .clk(b0mlcn000hn1n02x5_66_clk),
    .o(b0mlcn000hn1n02x5_66_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_67 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_67_d),
    .clk(b0mlcn000hn1n02x5_67_clk),
    .o(b0mlcn000hn1n02x5_67_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_68 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_68_d),
    .clk(b0mlcn000hn1n02x5_68_clk),
    .o(b0mlcn000hn1n02x5_68_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_69 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_69_d),
    .clk(b0mlcn000hn1n02x5_69_clk),
    .o(b0mlcn000hn1n02x5_69_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_70 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_70_d),
    .clk(b0mlcn000hn1n02x5_70_clk),
    .o(b0mlcn000hn1n02x5_70_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_71 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_71_d),
    .clk(b0mlcn000hn1n02x5_71_clk),
    .o(b0mlcn000hn1n02x5_71_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_72 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_72_d),
    .clk(b0mlcn000hn1n02x5_72_clk),
    .o(b0mlcn000hn1n02x5_72_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_73 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_73_d),
    .clk(b0mlcn000hn1n02x5_73_clk),
    .o(b0mlcn000hn1n02x5_73_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_74 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_74_d),
    .clk(b0mlcn000hn1n02x5_74_clk),
    .o(b0mlcn000hn1n02x5_74_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_75 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_75_d),
    .clk(b0mlcn000hn1n02x5_75_clk),
    .o(b0mlcn000hn1n02x5_75_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_76 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_76_d),
    .clk(b0mlcn000hn1n02x5_76_clk),
    .o(b0mlcn000hn1n02x5_76_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_77 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_77_d),
    .clk(b0mlcn000hn1n02x5_77_clk),
    .o(b0mlcn000hn1n02x5_77_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_78 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_78_d),
    .clk(b0mlcn000hn1n02x5_78_clk),
    .o(b0mlcn000hn1n02x5_78_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_79 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_79_d),
    .clk(b0mlcn000hn1n02x5_79_clk),
    .o(b0mlcn000hn1n02x5_79_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_80 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_80_d),
    .clk(b0mlcn000hn1n02x5_80_clk),
    .o(b0mlcn000hn1n02x5_80_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_81 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_81_d),
    .clk(b0mlcn000hn1n02x5_81_clk),
    .o(b0mlcn000hn1n02x5_81_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_82 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_82_d),
    .clk(b0mlcn000hn1n02x5_82_clk),
    .o(b0mlcn000hn1n02x5_82_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_83 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_83_d),
    .clk(b0mlcn000hn1n02x5_83_clk),
    .o(b0mlcn000hn1n02x5_83_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_84 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_84_d),
    .clk(b0mlcn000hn1n02x5_84_clk),
    .o(b0mlcn000hn1n02x5_84_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_85 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_85_d),
    .clk(b0mlcn000hn1n02x5_85_clk),
    .o(b0mlcn000hn1n02x5_85_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_86 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_86_d),
    .clk(b0mlcn000hn1n02x5_86_clk),
    .o(b0mlcn000hn1n02x5_86_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_87 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_87_d),
    .clk(b0mlcn000hn1n02x5_87_clk),
    .o(b0mlcn000hn1n02x5_87_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_88 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_88_d),
    .clk(b0mlcn000hn1n02x5_88_clk),
    .o(b0mlcn000hn1n02x5_88_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_89 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_89_d),
    .clk(b0mlcn000hn1n02x5_89_clk),
    .o(b0mlcn000hn1n02x5_89_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_90 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_90_d),
    .clk(b0mlcn000hn1n02x5_90_clk),
    .o(b0mlcn000hn1n02x5_90_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_91 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_91_d),
    .clk(b0mlcn000hn1n02x5_91_clk),
    .o(b0mlcn000hn1n02x5_91_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_92 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_92_d),
    .clk(b0mlcn000hn1n02x5_92_clk),
    .o(b0mlcn000hn1n02x5_92_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_93 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_93_d),
    .clk(b0mlcn000hn1n02x5_93_clk),
    .o(b0mlcn000hn1n02x5_93_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_94 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_94_d),
    .clk(b0mlcn000hn1n02x5_94_clk),
    .o(b0mlcn000hn1n02x5_94_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_95 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_95_d),
    .clk(b0mlcn000hn1n02x5_95_clk),
    .o(b0mlcn000hn1n02x5_95_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_96 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_96_d),
    .clk(b0mlcn000hn1n02x5_96_clk),
    .o(b0mlcn000hn1n02x5_96_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_97 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_97_d),
    .clk(b0mlcn000hn1n02x5_97_clk),
    .o(b0mlcn000hn1n02x5_97_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_98 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_98_d),
    .clk(b0mlcn000hn1n02x5_98_clk),
    .o(b0mlcn000hn1n02x5_98_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_99 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_99_d),
    .clk(b0mlcn000hn1n02x5_99_clk),
    .o(b0mlcn000hn1n02x5_99_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_100 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_100_d),
    .clk(b0mlcn000hn1n02x5_100_clk),
    .o(b0mlcn000hn1n02x5_100_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_101 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_101_d),
    .clk(b0mlcn000hn1n02x5_101_clk),
    .o(b0mlcn000hn1n02x5_101_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_102 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_102_d),
    .clk(b0mlcn000hn1n02x5_102_clk),
    .o(b0mlcn000hn1n02x5_102_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_103 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_103_d),
    .clk(b0mlcn000hn1n02x5_103_clk),
    .o(b0mlcn000hn1n02x5_103_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_104 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_104_d),
    .clk(b0mlcn000hn1n02x5_104_clk),
    .o(b0mlcn000hn1n02x5_104_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_105 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_105_d),
    .clk(b0mlcn000hn1n02x5_105_clk),
    .o(b0mlcn000hn1n02x5_105_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_106 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_106_d),
    .clk(b0mlcn000hn1n02x5_106_clk),
    .o(b0mlcn000hn1n02x5_106_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_107 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_107_d),
    .clk(b0mlcn000hn1n02x5_107_clk),
    .o(b0mlcn000hn1n02x5_107_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_108 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_108_d),
    .clk(b0mlcn000hn1n02x5_108_clk),
    .o(b0mlcn000hn1n02x5_108_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_109 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_109_d),
    .clk(b0mlcn000hn1n02x5_109_clk),
    .o(b0mlcn000hn1n02x5_109_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_110 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_110_d),
    .clk(b0mlcn000hn1n02x5_110_clk),
    .o(b0mlcn000hn1n02x5_110_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_111 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_111_d),
    .clk(b0mlcn000hn1n02x5_111_clk),
    .o(b0mlcn000hn1n02x5_111_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_112 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_112_d),
    .clk(b0mlcn000hn1n02x5_112_clk),
    .o(b0mlcn000hn1n02x5_112_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_113 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_113_d),
    .clk(b0mlcn000hn1n02x5_113_clk),
    .o(b0mlcn000hn1n02x5_113_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_114 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_114_d),
    .clk(b0mlcn000hn1n02x5_114_clk),
    .o(b0mlcn000hn1n02x5_114_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_115 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_115_d),
    .clk(b0mlcn000hn1n02x5_115_clk),
    .o(b0mlcn000hn1n02x5_115_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_116 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_116_d),
    .clk(b0mlcn000hn1n02x5_116_clk),
    .o(b0mlcn000hn1n02x5_116_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_117 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_117_d),
    .clk(b0mlcn000hn1n02x5_117_clk),
    .o(b0mlcn000hn1n02x5_117_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_118 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_118_d),
    .clk(b0mlcn000hn1n02x5_118_clk),
    .o(b0mlcn000hn1n02x5_118_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_119 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_119_d),
    .clk(b0mlcn000hn1n02x5_119_clk),
    .o(b0mlcn000hn1n02x5_119_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_120 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_120_d),
    .clk(b0mlcn000hn1n02x5_120_clk),
    .o(b0mlcn000hn1n02x5_120_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_121 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_121_d),
    .clk(b0mlcn000hn1n02x5_121_clk),
    .o(b0mlcn000hn1n02x5_121_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_122 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_122_d),
    .clk(b0mlcn000hn1n02x5_122_clk),
    .o(b0mlcn000hn1n02x5_122_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_123 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_123_d),
    .clk(b0mlcn000hn1n02x5_123_clk),
    .o(b0mlcn000hn1n02x5_123_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_124 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_124_d),
    .clk(b0mlcn000hn1n02x5_124_clk),
    .o(b0mlcn000hn1n02x5_124_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_125 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_125_d),
    .clk(b0mlcn000hn1n02x5_125_clk),
    .o(b0mlcn000hn1n02x5_125_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_126 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_126_d),
    .clk(b0mlcn000hn1n02x5_126_clk),
    .o(b0mlcn000hn1n02x5_126_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_127 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_127_d),
    .clk(b0mlcn000hn1n02x5_127_clk),
    .o(b0mlcn000hn1n02x5_127_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_128 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_128_d),
    .clk(b0mlcn000hn1n02x5_128_clk),
    .o(b0mlcn000hn1n02x5_128_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_129 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_129_d),
    .clk(b0mlcn000hn1n02x5_129_clk),
    .o(b0mlcn000hn1n02x5_129_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_130 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_130_d),
    .clk(b0mlcn000hn1n02x5_130_clk),
    .o(b0mlcn000hn1n02x5_130_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_131 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_131_d),
    .clk(b0mlcn000hn1n02x5_131_clk),
    .o(b0mlcn000hn1n02x5_131_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_132 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_132_d),
    .clk(b0mlcn000hn1n02x5_132_clk),
    .o(b0mlcn000hn1n02x5_132_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_133 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_133_d),
    .clk(b0mlcn000hn1n02x5_133_clk),
    .o(b0mlcn000hn1n02x5_133_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_134 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_134_d),
    .clk(b0mlcn000hn1n02x5_134_clk),
    .o(b0mlcn000hn1n02x5_134_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_135 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_135_d),
    .clk(b0mlcn000hn1n02x5_135_clk),
    .o(b0mlcn000hn1n02x5_135_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_136 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_136_d),
    .clk(b0mlcn000hn1n02x5_136_clk),
    .o(b0mlcn000hn1n02x5_136_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_137 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_137_d),
    .clk(b0mlcn000hn1n02x5_137_clk),
    .o(b0mlcn000hn1n02x5_137_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_138 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_138_d),
    .clk(b0mlcn000hn1n02x5_138_clk),
    .o(b0mlcn000hn1n02x5_138_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_139 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_139_d),
    .clk(b0mlcn000hn1n02x5_139_clk),
    .o(b0mlcn000hn1n02x5_139_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_140 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_140_d),
    .clk(b0mlcn000hn1n02x5_140_clk),
    .o(b0mlcn000hn1n02x5_140_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_141 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_141_d),
    .clk(b0mlcn000hn1n02x5_141_clk),
    .o(b0mlcn000hn1n02x5_141_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_142 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_142_d),
    .clk(b0mlcn000hn1n02x5_142_clk),
    .o(b0mlcn000hn1n02x5_142_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_143 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_143_d),
    .clk(b0mlcn000hn1n02x5_143_clk),
    .o(b0mlcn000hn1n02x5_143_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_144 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_144_d),
    .clk(b0mlcn000hn1n02x5_144_clk),
    .o(b0mlcn000hn1n02x5_144_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_145 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_145_d),
    .clk(b0mlcn000hn1n02x5_145_clk),
    .o(b0mlcn000hn1n02x5_145_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_146 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_146_d),
    .clk(b0mlcn000hn1n02x5_146_clk),
    .o(b0mlcn000hn1n02x5_146_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_147 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_147_d),
    .clk(b0mlcn000hn1n02x5_147_clk),
    .o(b0mlcn000hn1n02x5_147_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_148 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_148_d),
    .clk(b0mlcn000hn1n02x5_148_clk),
    .o(b0mlcn000hn1n02x5_148_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_149 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_149_d),
    .clk(b0mlcn000hn1n02x5_149_clk),
    .o(b0mlcn000hn1n02x5_149_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_150 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_150_d),
    .clk(b0mlcn000hn1n02x5_150_clk),
    .o(b0mlcn000hn1n02x5_150_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_151 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_151_d),
    .clk(b0mlcn000hn1n02x5_151_clk),
    .o(b0mlcn000hn1n02x5_151_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_152 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_152_d),
    .clk(b0mlcn000hn1n02x5_152_clk),
    .o(b0mlcn000hn1n02x5_152_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_153 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_153_d),
    .clk(b0mlcn000hn1n02x5_153_clk),
    .o(b0mlcn000hn1n02x5_153_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_154 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_154_d),
    .clk(b0mlcn000hn1n02x5_154_clk),
    .o(b0mlcn000hn1n02x5_154_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_155 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_155_d),
    .clk(b0mlcn000hn1n02x5_155_clk),
    .o(b0mlcn000hn1n02x5_155_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_156 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_156_d),
    .clk(b0mlcn000hn1n02x5_156_clk),
    .o(b0mlcn000hn1n02x5_156_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_157 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_157_d),
    .clk(b0mlcn000hn1n02x5_157_clk),
    .o(b0mlcn000hn1n02x5_157_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_158 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_158_d),
    .clk(b0mlcn000hn1n02x5_158_clk),
    .o(b0mlcn000hn1n02x5_158_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_159 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_159_d),
    .clk(b0mlcn000hn1n02x5_159_clk),
    .o(b0mlcn000hn1n02x5_159_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_160 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_160_d),
    .clk(b0mlcn000hn1n02x5_160_clk),
    .o(b0mlcn000hn1n02x5_160_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_161 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_161_d),
    .clk(b0mlcn000hn1n02x5_161_clk),
    .o(b0mlcn000hn1n02x5_161_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_162 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_162_d),
    .clk(b0mlcn000hn1n02x5_162_clk),
    .o(b0mlcn000hn1n02x5_162_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_163 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_163_d),
    .clk(b0mlcn000hn1n02x5_163_clk),
    .o(b0mlcn000hn1n02x5_163_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_164 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_164_d),
    .clk(b0mlcn000hn1n02x5_164_clk),
    .o(b0mlcn000hn1n02x5_164_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_165 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_165_d),
    .clk(b0mlcn000hn1n02x5_165_clk),
    .o(b0mlcn000hn1n02x5_165_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_166 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_166_d),
    .clk(b0mlcn000hn1n02x5_166_clk),
    .o(b0mlcn000hn1n02x5_166_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_167 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_167_d),
    .clk(b0mlcn000hn1n02x5_167_clk),
    .o(b0mlcn000hn1n02x5_167_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_168 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_168_d),
    .clk(b0mlcn000hn1n02x5_168_clk),
    .o(b0mlcn000hn1n02x5_168_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_169 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_169_d),
    .clk(b0mlcn000hn1n02x5_169_clk),
    .o(b0mlcn000hn1n02x5_169_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_170 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_170_d),
    .clk(b0mlcn000hn1n02x5_170_clk),
    .o(b0mlcn000hn1n02x5_170_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_171 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_171_d),
    .clk(b0mlcn000hn1n02x5_171_clk),
    .o(b0mlcn000hn1n02x5_171_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_172 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_172_d),
    .clk(b0mlcn000hn1n02x5_172_clk),
    .o(b0mlcn000hn1n02x5_172_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_173 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_173_d),
    .clk(b0mlcn000hn1n02x5_173_clk),
    .o(b0mlcn000hn1n02x5_173_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_174 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_174_d),
    .clk(b0mlcn000hn1n02x5_174_clk),
    .o(b0mlcn000hn1n02x5_174_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_175 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_175_d),
    .clk(b0mlcn000hn1n02x5_175_clk),
    .o(b0mlcn000hn1n02x5_175_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_176 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_176_d),
    .clk(b0mlcn000hn1n02x5_176_clk),
    .o(b0mlcn000hn1n02x5_176_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_177 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_177_d),
    .clk(b0mlcn000hn1n02x5_177_clk),
    .o(b0mlcn000hn1n02x5_177_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_178 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_178_d),
    .clk(b0mlcn000hn1n02x5_178_clk),
    .o(b0mlcn000hn1n02x5_178_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_179 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_179_d),
    .clk(b0mlcn000hn1n02x5_179_clk),
    .o(b0mlcn000hn1n02x5_179_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_180 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_180_d),
    .clk(b0mlcn000hn1n02x5_180_clk),
    .o(b0mlcn000hn1n02x5_180_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_181 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_181_d),
    .clk(b0mlcn000hn1n02x5_181_clk),
    .o(b0mlcn000hn1n02x5_181_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_182 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_182_d),
    .clk(b0mlcn000hn1n02x5_182_clk),
    .o(b0mlcn000hn1n02x5_182_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_183 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_183_d),
    .clk(b0mlcn000hn1n02x5_183_clk),
    .o(b0mlcn000hn1n02x5_183_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_184 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_184_d),
    .clk(b0mlcn000hn1n02x5_184_clk),
    .o(b0mlcn000hn1n02x5_184_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_185 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_185_d),
    .clk(b0mlcn000hn1n02x5_185_clk),
    .o(b0mlcn000hn1n02x5_185_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_186 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_186_d),
    .clk(b0mlcn000hn1n02x5_186_clk),
    .o(b0mlcn000hn1n02x5_186_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_187 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_187_d),
    .clk(b0mlcn000hn1n02x5_187_clk),
    .o(b0mlcn000hn1n02x5_187_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_188 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_188_d),
    .clk(b0mlcn000hn1n02x5_188_clk),
    .o(b0mlcn000hn1n02x5_188_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_189 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_189_d),
    .clk(b0mlcn000hn1n02x5_189_clk),
    .o(b0mlcn000hn1n02x5_189_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_190 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_190_d),
    .clk(b0mlcn000hn1n02x5_190_clk),
    .o(b0mlcn000hn1n02x5_190_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_191 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_191_d),
    .clk(b0mlcn000hn1n02x5_191_clk),
    .o(b0mlcn000hn1n02x5_191_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_192 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_192_d),
    .clk(b0mlcn000hn1n02x5_192_clk),
    .o(b0mlcn000hn1n02x5_192_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_193 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_193_d),
    .clk(b0mlcn000hn1n02x5_193_clk),
    .o(b0mlcn000hn1n02x5_193_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_194 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_194_d),
    .clk(b0mlcn000hn1n02x5_194_clk),
    .o(b0mlcn000hn1n02x5_194_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_195 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_195_d),
    .clk(b0mlcn000hn1n02x5_195_clk),
    .o(b0mlcn000hn1n02x5_195_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_196 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_196_d),
    .clk(b0mlcn000hn1n02x5_196_clk),
    .o(b0mlcn000hn1n02x5_196_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_197 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_197_d),
    .clk(b0mlcn000hn1n02x5_197_clk),
    .o(b0mlcn000hn1n02x5_197_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_198 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_198_d),
    .clk(b0mlcn000hn1n02x5_198_clk),
    .o(b0mlcn000hn1n02x5_198_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_199 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_199_d),
    .clk(b0mlcn000hn1n02x5_199_clk),
    .o(b0mlcn000hn1n02x5_199_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_200 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_200_d),
    .clk(b0mlcn000hn1n02x5_200_clk),
    .o(b0mlcn000hn1n02x5_200_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_201 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_201_d),
    .clk(b0mlcn000hn1n02x5_201_clk),
    .o(b0mlcn000hn1n02x5_201_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_202 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_202_d),
    .clk(b0mlcn000hn1n02x5_202_clk),
    .o(b0mlcn000hn1n02x5_202_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_203 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_203_d),
    .clk(b0mlcn000hn1n02x5_203_clk),
    .o(b0mlcn000hn1n02x5_203_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_204 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_204_d),
    .clk(b0mlcn000hn1n02x5_204_clk),
    .o(b0mlcn000hn1n02x5_204_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_205 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_205_d),
    .clk(b0mlcn000hn1n02x5_205_clk),
    .o(b0mlcn000hn1n02x5_205_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_206 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_206_d),
    .clk(b0mlcn000hn1n02x5_206_clk),
    .o(b0mlcn000hn1n02x5_206_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_207 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_207_d),
    .clk(b0mlcn000hn1n02x5_207_clk),
    .o(b0mlcn000hn1n02x5_207_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_208 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_208_d),
    .clk(b0mlcn000hn1n02x5_208_clk),
    .o(b0mlcn000hn1n02x5_208_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_209 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_209_d),
    .clk(b0mlcn000hn1n02x5_209_clk),
    .o(b0mlcn000hn1n02x5_209_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_210 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_210_d),
    .clk(b0mlcn000hn1n02x5_210_clk),
    .o(b0mlcn000hn1n02x5_210_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_211 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_211_d),
    .clk(b0mlcn000hn1n02x5_211_clk),
    .o(b0mlcn000hn1n02x5_211_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_212 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_212_d),
    .clk(b0mlcn000hn1n02x5_212_clk),
    .o(b0mlcn000hn1n02x5_212_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_213 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_213_d),
    .clk(b0mlcn000hn1n02x5_213_clk),
    .o(b0mlcn000hn1n02x5_213_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_214 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_214_d),
    .clk(b0mlcn000hn1n02x5_214_clk),
    .o(b0mlcn000hn1n02x5_214_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_215 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_215_d),
    .clk(b0mlcn000hn1n02x5_215_clk),
    .o(b0mlcn000hn1n02x5_215_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_216 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_216_d),
    .clk(b0mlcn000hn1n02x5_216_clk),
    .o(b0mlcn000hn1n02x5_216_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_217 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_217_d),
    .clk(b0mlcn000hn1n02x5_217_clk),
    .o(b0mlcn000hn1n02x5_217_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_218 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_218_d),
    .clk(b0mlcn000hn1n02x5_218_clk),
    .o(b0mlcn000hn1n02x5_218_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_219 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_219_d),
    .clk(b0mlcn000hn1n02x5_219_clk),
    .o(b0mlcn000hn1n02x5_219_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_220 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_220_d),
    .clk(b0mlcn000hn1n02x5_220_clk),
    .o(b0mlcn000hn1n02x5_220_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_221 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_221_d),
    .clk(b0mlcn000hn1n02x5_221_clk),
    .o(b0mlcn000hn1n02x5_221_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_222 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_222_d),
    .clk(b0mlcn000hn1n02x5_222_clk),
    .o(b0mlcn000hn1n02x5_222_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_223 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_223_d),
    .clk(b0mlcn000hn1n02x5_223_clk),
    .o(b0mlcn000hn1n02x5_223_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_224 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_224_d),
    .clk(b0mlcn000hn1n02x5_224_clk),
    .o(b0mlcn000hn1n02x5_224_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_225 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_225_d),
    .clk(b0mlcn000hn1n02x5_225_clk),
    .o(b0mlcn000hn1n02x5_225_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_226 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_226_d),
    .clk(b0mlcn000hn1n02x5_226_clk),
    .o(b0mlcn000hn1n02x5_226_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_227 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_227_d),
    .clk(b0mlcn000hn1n02x5_227_clk),
    .o(b0mlcn000hn1n02x5_227_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_228 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_228_d),
    .clk(b0mlcn000hn1n02x5_228_clk),
    .o(b0mlcn000hn1n02x5_228_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_229 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_229_d),
    .clk(b0mlcn000hn1n02x5_229_clk),
    .o(b0mlcn000hn1n02x5_229_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_230 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_230_d),
    .clk(b0mlcn000hn1n02x5_230_clk),
    .o(b0mlcn000hn1n02x5_230_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_231 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_231_d),
    .clk(b0mlcn000hn1n02x5_231_clk),
    .o(b0mlcn000hn1n02x5_231_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_232 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_232_d),
    .clk(b0mlcn000hn1n02x5_232_clk),
    .o(b0mlcn000hn1n02x5_232_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_233 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_233_d),
    .clk(b0mlcn000hn1n02x5_233_clk),
    .o(b0mlcn000hn1n02x5_233_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_234 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_234_d),
    .clk(b0mlcn000hn1n02x5_234_clk),
    .o(b0mlcn000hn1n02x5_234_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_235 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_235_d),
    .clk(b0mlcn000hn1n02x5_235_clk),
    .o(b0mlcn000hn1n02x5_235_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_236 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_236_d),
    .clk(b0mlcn000hn1n02x5_236_clk),
    .o(b0mlcn000hn1n02x5_236_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_237 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_237_d),
    .clk(b0mlcn000hn1n02x5_237_clk),
    .o(b0mlcn000hn1n02x5_237_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_238 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_238_d),
    .clk(b0mlcn000hn1n02x5_238_clk),
    .o(b0mlcn000hn1n02x5_238_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_239 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_239_d),
    .clk(b0mlcn000hn1n02x5_239_clk),
    .o(b0mlcn000hn1n02x5_239_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_240 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_240_d),
    .clk(b0mlcn000hn1n02x5_240_clk),
    .o(b0mlcn000hn1n02x5_240_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_241 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_241_d),
    .clk(b0mlcn000hn1n02x5_241_clk),
    .o(b0mlcn000hn1n02x5_241_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_242 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_242_d),
    .clk(b0mlcn000hn1n02x5_242_clk),
    .o(b0mlcn000hn1n02x5_242_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_243 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_243_d),
    .clk(b0mlcn000hn1n02x5_243_clk),
    .o(b0mlcn000hn1n02x5_243_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_244 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_244_d),
    .clk(b0mlcn000hn1n02x5_244_clk),
    .o(b0mlcn000hn1n02x5_244_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_245 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_245_d),
    .clk(b0mlcn000hn1n02x5_245_clk),
    .o(b0mlcn000hn1n02x5_245_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_246 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_246_d),
    .clk(b0mlcn000hn1n02x5_246_clk),
    .o(b0mlcn000hn1n02x5_246_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_247 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_247_d),
    .clk(b0mlcn000hn1n02x5_247_clk),
    .o(b0mlcn000hn1n02x5_247_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_248 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_248_d),
    .clk(b0mlcn000hn1n02x5_248_clk),
    .o(b0mlcn000hn1n02x5_248_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_249 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_249_d),
    .clk(b0mlcn000hn1n02x5_249_clk),
    .o(b0mlcn000hn1n02x5_249_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_250 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_250_d),
    .clk(b0mlcn000hn1n02x5_250_clk),
    .o(b0mlcn000hn1n02x5_250_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_251 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_251_d),
    .clk(b0mlcn000hn1n02x5_251_clk),
    .o(b0mlcn000hn1n02x5_251_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_252 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_252_d),
    .clk(b0mlcn000hn1n02x5_252_clk),
    .o(b0mlcn000hn1n02x5_252_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_253 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_253_d),
    .clk(b0mlcn000hn1n02x5_253_clk),
    .o(b0mlcn000hn1n02x5_253_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_254 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_254_d),
    .clk(b0mlcn000hn1n02x5_254_clk),
    .o(b0mlcn000hn1n02x5_254_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_255 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_255_d),
    .clk(b0mlcn000hn1n02x5_255_clk),
    .o(b0mlcn000hn1n02x5_255_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_256 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_256_d),
    .clk(b0mlcn000hn1n02x5_256_clk),
    .o(b0mlcn000hn1n02x5_256_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_257 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_257_d),
    .clk(b0mlcn000hn1n02x5_257_clk),
    .o(b0mlcn000hn1n02x5_257_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_258 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_258_d),
    .clk(b0mlcn000hn1n02x5_258_clk),
    .o(b0mlcn000hn1n02x5_258_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_259 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_259_d),
    .clk(b0mlcn000hn1n02x5_259_clk),
    .o(b0mlcn000hn1n02x5_259_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_260 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_260_d),
    .clk(b0mlcn000hn1n02x5_260_clk),
    .o(b0mlcn000hn1n02x5_260_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_261 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_261_d),
    .clk(b0mlcn000hn1n02x5_261_clk),
    .o(b0mlcn000hn1n02x5_261_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_262 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_262_d),
    .clk(b0mlcn000hn1n02x5_262_clk),
    .o(b0mlcn000hn1n02x5_262_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_263 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_263_d),
    .clk(b0mlcn000hn1n02x5_263_clk),
    .o(b0mlcn000hn1n02x5_263_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_264 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_264_d),
    .clk(b0mlcn000hn1n02x5_264_clk),
    .o(b0mlcn000hn1n02x5_264_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_265 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_265_d),
    .clk(b0mlcn000hn1n02x5_265_clk),
    .o(b0mlcn000hn1n02x5_265_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_266 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_266_d),
    .clk(b0mlcn000hn1n02x5_266_clk),
    .o(b0mlcn000hn1n02x5_266_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_267 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_267_d),
    .clk(b0mlcn000hn1n02x5_267_clk),
    .o(b0mlcn000hn1n02x5_267_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_268 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_268_d),
    .clk(b0mlcn000hn1n02x5_268_clk),
    .o(b0mlcn000hn1n02x5_268_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_269 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_269_d),
    .clk(b0mlcn000hn1n02x5_269_clk),
    .o(b0mlcn000hn1n02x5_269_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_270 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_270_d),
    .clk(b0mlcn000hn1n02x5_270_clk),
    .o(b0mlcn000hn1n02x5_270_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_271 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_271_d),
    .clk(b0mlcn000hn1n02x5_271_clk),
    .o(b0mlcn000hn1n02x5_271_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_272 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_272_d),
    .clk(b0mlcn000hn1n02x5_272_clk),
    .o(b0mlcn000hn1n02x5_272_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_273 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_273_d),
    .clk(b0mlcn000hn1n02x5_273_clk),
    .o(b0mlcn000hn1n02x5_273_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_274 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_274_d),
    .clk(b0mlcn000hn1n02x5_274_clk),
    .o(b0mlcn000hn1n02x5_274_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_275 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_275_d),
    .clk(b0mlcn000hn1n02x5_275_clk),
    .o(b0mlcn000hn1n02x5_275_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_276 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_276_d),
    .clk(b0mlcn000hn1n02x5_276_clk),
    .o(b0mlcn000hn1n02x5_276_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_277 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_277_d),
    .clk(b0mlcn000hn1n02x5_277_clk),
    .o(b0mlcn000hn1n02x5_277_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_278 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_278_d),
    .clk(b0mlcn000hn1n02x5_278_clk),
    .o(b0mlcn000hn1n02x5_278_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_279 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_279_d),
    .clk(b0mlcn000hn1n02x5_279_clk),
    .o(b0mlcn000hn1n02x5_279_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_280 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_280_d),
    .clk(b0mlcn000hn1n02x5_280_clk),
    .o(b0mlcn000hn1n02x5_280_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_281 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_281_d),
    .clk(b0mlcn000hn1n02x5_281_clk),
    .o(b0mlcn000hn1n02x5_281_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_282 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_282_d),
    .clk(b0mlcn000hn1n02x5_282_clk),
    .o(b0mlcn000hn1n02x5_282_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_283 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_283_d),
    .clk(b0mlcn000hn1n02x5_283_clk),
    .o(b0mlcn000hn1n02x5_283_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_284 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_284_d),
    .clk(b0mlcn000hn1n02x5_284_clk),
    .o(b0mlcn000hn1n02x5_284_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_285 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_285_d),
    .clk(b0mlcn000hn1n02x5_285_clk),
    .o(b0mlcn000hn1n02x5_285_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_286 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_286_d),
    .clk(b0mlcn000hn1n02x5_286_clk),
    .o(b0mlcn000hn1n02x5_286_o)
  );
  b0mlcn000hn1n02x5 b0mlcn000hn1n02x5_287 ( // @[ScanConfRadh.scala 61:46]
    .d(b0mlcn000hn1n02x5_287_d),
    .clk(b0mlcn000hn1n02x5_287_clk),
    .o(b0mlcn000hn1n02x5_287_o)
  );
  assign ioBundle_confOut = {io_confOut_hi,io_confOut_lo}; // @[ScanConfRadh.scala 67:45]
  assign ioBundle_scan_out = {io_scan_out_hi,io_scan_out_lo}; // @[ScanConfRadh.scala 59:47]
  assign b0mlcn000hn1n02x5_d = confReg_0; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_1_d = confReg_1; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_1_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_2_d = confReg_2; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_2_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_3_d = confReg_3; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_3_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_4_d = confReg_4; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_4_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_5_d = confReg_5; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_5_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_6_d = confReg_6; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_6_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_7_d = confReg_7; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_7_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_8_d = confReg_8; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_8_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_9_d = confReg_9; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_9_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_10_d = confReg_10; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_10_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_11_d = confReg_11; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_11_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_12_d = confReg_12; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_12_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_13_d = confReg_13; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_13_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_14_d = confReg_14; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_14_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_15_d = confReg_15; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_15_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_16_d = confReg_16; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_16_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_17_d = confReg_17; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_17_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_18_d = confReg_18; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_18_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_19_d = confReg_19; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_19_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_20_d = confReg_20; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_20_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_21_d = confReg_21; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_21_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_22_d = confReg_22; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_22_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_23_d = confReg_23; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_23_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_24_d = confReg_24; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_24_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_25_d = confReg_25; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_25_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_26_d = confReg_26; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_26_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_27_d = confReg_27; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_27_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_28_d = confReg_28; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_28_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_29_d = confReg_29; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_29_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_30_d = confReg_30; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_30_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_31_d = confReg_31; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_31_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_32_d = confReg_32; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_32_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_33_d = confReg_33; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_33_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_34_d = confReg_34; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_34_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_35_d = confReg_35; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_35_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_36_d = confReg_36; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_36_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_37_d = confReg_37; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_37_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_38_d = confReg_38; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_38_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_39_d = confReg_39; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_39_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_40_d = confReg_40; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_40_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_41_d = confReg_41; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_41_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_42_d = confReg_42; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_42_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_43_d = confReg_43; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_43_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_44_d = confReg_44; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_44_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_45_d = confReg_45; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_45_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_46_d = confReg_46; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_46_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_47_d = confReg_47; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_47_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_48_d = confReg_48; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_48_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_49_d = confReg_49; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_49_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_50_d = confReg_50; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_50_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_51_d = confReg_51; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_51_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_52_d = confReg_52; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_52_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_53_d = confReg_53; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_53_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_54_d = confReg_54; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_54_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_55_d = confReg_55; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_55_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_56_d = confReg_56; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_56_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_57_d = confReg_57; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_57_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_58_d = confReg_58; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_58_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_59_d = confReg_59; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_59_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_60_d = confReg_60; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_60_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_61_d = confReg_61; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_61_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_62_d = confReg_62; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_62_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_63_d = confReg_63; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_63_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_64_d = confReg_64; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_64_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_65_d = confReg_65; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_65_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_66_d = confReg_66; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_66_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_67_d = confReg_67; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_67_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_68_d = confReg_68; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_68_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_69_d = confReg_69; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_69_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_70_d = confReg_70; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_70_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_71_d = confReg_71; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_71_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_72_d = confReg_72; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_72_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_73_d = confReg_73; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_73_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_74_d = confReg_74; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_74_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_75_d = confReg_75; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_75_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_76_d = confReg_76; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_76_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_77_d = confReg_77; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_77_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_78_d = confReg_78; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_78_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_79_d = confReg_79; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_79_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_80_d = confReg_80; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_80_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_81_d = confReg_81; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_81_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_82_d = confReg_82; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_82_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_83_d = confReg_83; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_83_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_84_d = confReg_84; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_84_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_85_d = confReg_85; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_85_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_86_d = confReg_86; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_86_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_87_d = confReg_87; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_87_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_88_d = confReg_88; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_88_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_89_d = confReg_89; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_89_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_90_d = confReg_90; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_90_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_91_d = confReg_91; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_91_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_92_d = confReg_92; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_92_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_93_d = confReg_93; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_93_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_94_d = confReg_94; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_94_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_95_d = confReg_95; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_95_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_96_d = confReg_96; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_96_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_97_d = confReg_97; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_97_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_98_d = confReg_98; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_98_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_99_d = confReg_99; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_99_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_100_d = confReg_100; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_100_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_101_d = confReg_101; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_101_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_102_d = confReg_102; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_102_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_103_d = confReg_103; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_103_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_104_d = confReg_104; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_104_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_105_d = confReg_105; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_105_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_106_d = confReg_106; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_106_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_107_d = confReg_107; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_107_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_108_d = confReg_108; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_108_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_109_d = confReg_109; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_109_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_110_d = confReg_110; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_110_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_111_d = confReg_111; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_111_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_112_d = confReg_112; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_112_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_113_d = confReg_113; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_113_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_114_d = confReg_114; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_114_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_115_d = confReg_115; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_115_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_116_d = confReg_116; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_116_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_117_d = confReg_117; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_117_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_118_d = confReg_118; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_118_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_119_d = confReg_119; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_119_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_120_d = confReg_120; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_120_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_121_d = confReg_121; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_121_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_122_d = confReg_122; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_122_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_123_d = confReg_123; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_123_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_124_d = confReg_124; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_124_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_125_d = confReg_125; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_125_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_126_d = confReg_126; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_126_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_127_d = confReg_127; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_127_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_128_d = confReg_128; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_128_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_129_d = confReg_129; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_129_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_130_d = confReg_130; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_130_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_131_d = confReg_131; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_131_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_132_d = confReg_132; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_132_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_133_d = confReg_133; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_133_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_134_d = confReg_134; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_134_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_135_d = confReg_135; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_135_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_136_d = confReg_136; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_136_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_137_d = confReg_137; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_137_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_138_d = confReg_138; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_138_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_139_d = confReg_139; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_139_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_140_d = confReg_140; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_140_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_141_d = confReg_141; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_141_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_142_d = confReg_142; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_142_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_143_d = confReg_143; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_143_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_144_d = confReg_144; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_144_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_145_d = confReg_145; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_145_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_146_d = confReg_146; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_146_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_147_d = confReg_147; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_147_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_148_d = confReg_148; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_148_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_149_d = confReg_149; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_149_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_150_d = confReg_150; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_150_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_151_d = confReg_151; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_151_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_152_d = confReg_152; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_152_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_153_d = confReg_153; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_153_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_154_d = confReg_154; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_154_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_155_d = confReg_155; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_155_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_156_d = confReg_156; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_156_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_157_d = confReg_157; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_157_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_158_d = confReg_158; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_158_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_159_d = confReg_159; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_159_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_160_d = confReg_160; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_160_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_161_d = confReg_161; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_161_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_162_d = confReg_162; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_162_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_163_d = confReg_163; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_163_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_164_d = confReg_164; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_164_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_165_d = confReg_165; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_165_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_166_d = confReg_166; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_166_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_167_d = confReg_167; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_167_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_168_d = confReg_168; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_168_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_169_d = confReg_169; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_169_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_170_d = confReg_170; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_170_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_171_d = confReg_171; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_171_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_172_d = confReg_172; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_172_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_173_d = confReg_173; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_173_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_174_d = confReg_174; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_174_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_175_d = confReg_175; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_175_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_176_d = confReg_176; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_176_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_177_d = confReg_177; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_177_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_178_d = confReg_178; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_178_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_179_d = confReg_179; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_179_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_180_d = confReg_180; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_180_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_181_d = confReg_181; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_181_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_182_d = confReg_182; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_182_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_183_d = confReg_183; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_183_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_184_d = confReg_184; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_184_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_185_d = confReg_185; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_185_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_186_d = confReg_186; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_186_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_187_d = confReg_187; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_187_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_188_d = confReg_188; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_188_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_189_d = confReg_189; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_189_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_190_d = confReg_190; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_190_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_191_d = confReg_191; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_191_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_192_d = confReg_192; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_192_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_193_d = confReg_193; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_193_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_194_d = confReg_194; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_194_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_195_d = confReg_195; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_195_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_196_d = confReg_196; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_196_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_197_d = confReg_197; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_197_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_198_d = confReg_198; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_198_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_199_d = confReg_199; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_199_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_200_d = confReg_200; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_200_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_201_d = confReg_201; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_201_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_202_d = confReg_202; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_202_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_203_d = confReg_203; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_203_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_204_d = confReg_204; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_204_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_205_d = confReg_205; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_205_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_206_d = confReg_206; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_206_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_207_d = confReg_207; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_207_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_208_d = confReg_208; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_208_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_209_d = confReg_209; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_209_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_210_d = confReg_210; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_210_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_211_d = confReg_211; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_211_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_212_d = confReg_212; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_212_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_213_d = confReg_213; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_213_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_214_d = confReg_214; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_214_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_215_d = confReg_215; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_215_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_216_d = confReg_216; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_216_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_217_d = confReg_217; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_217_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_218_d = confReg_218; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_218_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_219_d = confReg_219; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_219_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_220_d = confReg_220; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_220_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_221_d = confReg_221; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_221_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_222_d = confReg_222; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_222_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_223_d = confReg_223; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_223_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_224_d = confReg_224; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_224_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_225_d = confReg_225; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_225_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_226_d = confReg_226; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_226_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_227_d = confReg_227; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_227_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_228_d = confReg_228; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_228_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_229_d = confReg_229; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_229_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_230_d = confReg_230; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_230_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_231_d = confReg_231; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_231_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_232_d = confReg_232; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_232_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_233_d = confReg_233; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_233_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_234_d = confReg_234; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_234_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_235_d = confReg_235; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_235_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_236_d = confReg_236; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_236_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_237_d = confReg_237; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_237_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_238_d = confReg_238; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_238_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_239_d = confReg_239; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_239_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_240_d = confReg_240; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_240_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_241_d = confReg_241; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_241_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_242_d = confReg_242; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_242_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_243_d = confReg_243; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_243_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_244_d = confReg_244; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_244_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_245_d = confReg_245; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_245_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_246_d = confReg_246; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_246_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_247_d = confReg_247; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_247_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_248_d = confReg_248; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_248_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_249_d = confReg_249; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_249_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_250_d = confReg_250; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_250_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_251_d = confReg_251; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_251_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_252_d = confReg_252; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_252_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_253_d = confReg_253; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_253_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_254_d = confReg_254; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_254_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_255_d = confReg_255; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_255_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_256_d = confReg_256; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_256_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_257_d = confReg_257; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_257_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_258_d = confReg_258; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_258_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_259_d = confReg_259; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_259_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_260_d = confReg_260; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_260_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_261_d = confReg_261; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_261_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_262_d = confReg_262; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_262_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_263_d = confReg_263; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_263_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_264_d = confReg_264; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_264_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_265_d = confReg_265; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_265_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_266_d = confReg_266; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_266_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_267_d = confReg_267; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_267_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_268_d = confReg_268; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_268_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_269_d = confReg_269; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_269_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_270_d = confReg_270; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_270_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_271_d = confReg_271; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_271_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_272_d = confReg_272; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_272_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_273_d = confReg_273; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_273_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_274_d = confReg_274; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_274_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_275_d = confReg_275; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_275_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_276_d = confReg_276; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_276_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_277_d = confReg_277; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_277_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_278_d = confReg_278; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_278_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_279_d = confReg_279; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_279_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_280_d = confReg_280; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_280_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_281_d = confReg_281; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_281_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_282_d = confReg_282; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_282_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_283_d = confReg_283; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_283_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_284_d = confReg_284; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_284_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_285_d = confReg_285; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_285_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_286_d = confReg_286; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_286_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  assign b0mlcn000hn1n02x5_287_d = confReg_287; // @[ScanConfRadh.scala 65:22]
  assign b0mlcn000hn1n02x5_287_clk = ioBundle_scan_ioLatchEnb; // @[ScanConfRadh.scala 64:46]
  always @(posedge clock) begin
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_0 <= confReg_16; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_1 <= confReg_17; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_2 <= confReg_18; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_3 <= confReg_19; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_4 <= confReg_20; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_5 <= confReg_21; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_6 <= confReg_22; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_7 <= confReg_23; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_8 <= confReg_24; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_9 <= confReg_25; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_10 <= confReg_26; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_11 <= confReg_27; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_12 <= confReg_28; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_13 <= confReg_29; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_14 <= confReg_30; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_15 <= confReg_31; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_16 <= confReg_32; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_17 <= confReg_33; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_18 <= confReg_34; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_19 <= confReg_35; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_20 <= confReg_36; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_21 <= confReg_37; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_22 <= confReg_38; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_23 <= confReg_39; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_24 <= confReg_40; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_25 <= confReg_41; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_26 <= confReg_42; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_27 <= confReg_43; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_28 <= confReg_44; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_29 <= confReg_45; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_30 <= confReg_46; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_31 <= confReg_47; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_32 <= confReg_48; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_33 <= confReg_49; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_34 <= confReg_50; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_35 <= confReg_51; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_36 <= confReg_52; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_37 <= confReg_53; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_38 <= confReg_54; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_39 <= confReg_55; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_40 <= confReg_56; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_41 <= confReg_57; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_42 <= confReg_58; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_43 <= confReg_59; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_44 <= confReg_60; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_45 <= confReg_61; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_46 <= confReg_62; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_47 <= confReg_63; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_48 <= confReg_64; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_49 <= confReg_65; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_50 <= confReg_66; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_51 <= confReg_67; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_52 <= confReg_68; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_53 <= confReg_69; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_54 <= confReg_70; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_55 <= confReg_71; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_56 <= confReg_72; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_57 <= confReg_73; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_58 <= confReg_74; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_59 <= confReg_75; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_60 <= confReg_76; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_61 <= confReg_77; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_62 <= confReg_78; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_63 <= confReg_79; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_64 <= confReg_80; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_65 <= confReg_81; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_66 <= confReg_82; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_67 <= confReg_83; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_68 <= confReg_84; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_69 <= confReg_85; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_70 <= confReg_86; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_71 <= confReg_87; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_72 <= confReg_88; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_73 <= confReg_89; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_74 <= confReg_90; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_75 <= confReg_91; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_76 <= confReg_92; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_77 <= confReg_93; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_78 <= confReg_94; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_79 <= confReg_95; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_80 <= confReg_96; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_81 <= confReg_97; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_82 <= confReg_98; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_83 <= confReg_99; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_84 <= confReg_100; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_85 <= confReg_101; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_86 <= confReg_102; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_87 <= confReg_103; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_88 <= confReg_104; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_89 <= confReg_105; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_90 <= confReg_106; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_91 <= confReg_107; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_92 <= confReg_108; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_93 <= confReg_109; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_94 <= confReg_110; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_95 <= confReg_111; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_96 <= confReg_112; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_97 <= confReg_113; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_98 <= confReg_114; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_99 <= confReg_115; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_100 <= confReg_116; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_101 <= confReg_117; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_102 <= confReg_118; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_103 <= confReg_119; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_104 <= confReg_120; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_105 <= confReg_121; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_106 <= confReg_122; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_107 <= confReg_123; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_108 <= confReg_124; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_109 <= confReg_125; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_110 <= confReg_126; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_111 <= confReg_127; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_112 <= confReg_128; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_113 <= confReg_129; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_114 <= confReg_130; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_115 <= confReg_131; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_116 <= confReg_132; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_117 <= confReg_133; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_118 <= confReg_134; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_119 <= confReg_135; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_120 <= confReg_136; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_121 <= confReg_137; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_122 <= confReg_138; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_123 <= confReg_139; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_124 <= confReg_140; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_125 <= confReg_141; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_126 <= confReg_142; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_127 <= confReg_143; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_128 <= confReg_144; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_129 <= confReg_145; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_130 <= confReg_146; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_131 <= confReg_147; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_132 <= confReg_148; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_133 <= confReg_149; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_134 <= confReg_150; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_135 <= confReg_151; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_136 <= confReg_152; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_137 <= confReg_153; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_138 <= confReg_154; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_139 <= confReg_155; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_140 <= confReg_156; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_141 <= confReg_157; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_142 <= confReg_158; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_143 <= confReg_159; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_144 <= confReg_160; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_145 <= confReg_161; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_146 <= confReg_162; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_147 <= confReg_163; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_148 <= confReg_164; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_149 <= confReg_165; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_150 <= confReg_166; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_151 <= confReg_167; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_152 <= confReg_168; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_153 <= confReg_169; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_154 <= confReg_170; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_155 <= confReg_171; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_156 <= confReg_172; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_157 <= confReg_173; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_158 <= confReg_174; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_159 <= confReg_175; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_160 <= confReg_176; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_161 <= confReg_177; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_162 <= confReg_178; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_163 <= confReg_179; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_164 <= confReg_180; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_165 <= confReg_181; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_166 <= confReg_182; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_167 <= confReg_183; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_168 <= confReg_184; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_169 <= confReg_185; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_170 <= confReg_186; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_171 <= confReg_187; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_172 <= confReg_188; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_173 <= confReg_189; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_174 <= confReg_190; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_175 <= confReg_191; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_176 <= confReg_192; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_177 <= confReg_193; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_178 <= confReg_194; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_179 <= confReg_195; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_180 <= confReg_196; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_181 <= confReg_197; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_182 <= confReg_198; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_183 <= confReg_199; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_184 <= confReg_200; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_185 <= confReg_201; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_186 <= confReg_202; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_187 <= confReg_203; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_188 <= confReg_204; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_189 <= confReg_205; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_190 <= confReg_206; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_191 <= confReg_207; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_192 <= confReg_208; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_193 <= confReg_209; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_194 <= confReg_210; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_195 <= confReg_211; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_196 <= confReg_212; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_197 <= confReg_213; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_198 <= confReg_214; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_199 <= confReg_215; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_200 <= confReg_216; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_201 <= confReg_217; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_202 <= confReg_218; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_203 <= confReg_219; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_204 <= confReg_220; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_205 <= confReg_221; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_206 <= confReg_222; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_207 <= confReg_223; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_208 <= confReg_224; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_209 <= confReg_225; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_210 <= confReg_226; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_211 <= confReg_227; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_212 <= confReg_228; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_213 <= confReg_229; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_214 <= confReg_230; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_215 <= confReg_231; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_216 <= confReg_232; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_217 <= confReg_233; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_218 <= confReg_234; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_219 <= confReg_235; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_220 <= confReg_236; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_221 <= confReg_237; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_222 <= confReg_238; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_223 <= confReg_239; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_224 <= confReg_240; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_225 <= confReg_241; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_226 <= confReg_242; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_227 <= confReg_243; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_228 <= confReg_244; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_229 <= confReg_245; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_230 <= confReg_246; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_231 <= confReg_247; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_232 <= confReg_248; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_233 <= confReg_249; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_234 <= confReg_250; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_235 <= confReg_251; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_236 <= confReg_252; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_237 <= confReg_253; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_238 <= confReg_254; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_239 <= confReg_255; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_240 <= confReg_256; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_241 <= confReg_257; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_242 <= confReg_258; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_243 <= confReg_259; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_244 <= confReg_260; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_245 <= confReg_261; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_246 <= confReg_262; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_247 <= confReg_263; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_248 <= confReg_264; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_249 <= confReg_265; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_250 <= confReg_266; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_251 <= confReg_267; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_252 <= confReg_268; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_253 <= confReg_269; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_254 <= confReg_270; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_255 <= confReg_271; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_256 <= confReg_272; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_257 <= confReg_273; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_258 <= confReg_274; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_259 <= confReg_275; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_260 <= confReg_276; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_261 <= confReg_277; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_262 <= confReg_278; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_263 <= confReg_279; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_264 <= confReg_280; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_265 <= confReg_281; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_266 <= confReg_282; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_267 <= confReg_283; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_268 <= confReg_284; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_269 <= confReg_285; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_270 <= confReg_286; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_271 <= confReg_287; // @[ScanConfRadh.scala 54:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_272 <= ioBundle_scan_in[0]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_273 <= ioBundle_scan_in[1]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_274 <= ioBundle_scan_in[2]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_275 <= ioBundle_scan_in[3]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_276 <= ioBundle_scan_in[4]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_277 <= ioBundle_scan_in[5]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_278 <= ioBundle_scan_in[6]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_279 <= ioBundle_scan_in[7]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_280 <= ioBundle_scan_in[8]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_281 <= ioBundle_scan_in[9]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_282 <= ioBundle_scan_in[10]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_283 <= ioBundle_scan_in[11]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_284 <= ioBundle_scan_in[12]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_285 <= ioBundle_scan_in[13]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_286 <= ioBundle_scan_in[14]; // @[ScanConfRadh.scala 51:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConfRadh.scala 50:20]
      confReg_287 <= ioBundle_scan_in[15]; // @[ScanConfRadh.scala 51:72]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  confReg_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  confReg_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  confReg_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  confReg_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  confReg_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  confReg_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  confReg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  confReg_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  confReg_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  confReg_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  confReg_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  confReg_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  confReg_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  confReg_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  confReg_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  confReg_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  confReg_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  confReg_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  confReg_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  confReg_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  confReg_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  confReg_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  confReg_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  confReg_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  confReg_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  confReg_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  confReg_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  confReg_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  confReg_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  confReg_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  confReg_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  confReg_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  confReg_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  confReg_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  confReg_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  confReg_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  confReg_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  confReg_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  confReg_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  confReg_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  confReg_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  confReg_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  confReg_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  confReg_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  confReg_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  confReg_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  confReg_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  confReg_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  confReg_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  confReg_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  confReg_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  confReg_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  confReg_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  confReg_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  confReg_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  confReg_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  confReg_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  confReg_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  confReg_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  confReg_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  confReg_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  confReg_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  confReg_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  confReg_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  confReg_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  confReg_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  confReg_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  confReg_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  confReg_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  confReg_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  confReg_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  confReg_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  confReg_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  confReg_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  confReg_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  confReg_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  confReg_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  confReg_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  confReg_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  confReg_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  confReg_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  confReg_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  confReg_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  confReg_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  confReg_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  confReg_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  confReg_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  confReg_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  confReg_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  confReg_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  confReg_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  confReg_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  confReg_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  confReg_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  confReg_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  confReg_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  confReg_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  confReg_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  confReg_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  confReg_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  confReg_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  confReg_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  confReg_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  confReg_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  confReg_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  confReg_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  confReg_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  confReg_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  confReg_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  confReg_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  confReg_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  confReg_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  confReg_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  confReg_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  confReg_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  confReg_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  confReg_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  confReg_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  confReg_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  confReg_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  confReg_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  confReg_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  confReg_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  confReg_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  confReg_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  confReg_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  confReg_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  confReg_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  confReg_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  confReg_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  confReg_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  confReg_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  confReg_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  confReg_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  confReg_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  confReg_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  confReg_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  confReg_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  confReg_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  confReg_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  confReg_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  confReg_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  confReg_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  confReg_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  confReg_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  confReg_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  confReg_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  confReg_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  confReg_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  confReg_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  confReg_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  confReg_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  confReg_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  confReg_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  confReg_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  confReg_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  confReg_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  confReg_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  confReg_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  confReg_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  confReg_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  confReg_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  confReg_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  confReg_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  confReg_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  confReg_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  confReg_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  confReg_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  confReg_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  confReg_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  confReg_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  confReg_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  confReg_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  confReg_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  confReg_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  confReg_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  confReg_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  confReg_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  confReg_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  confReg_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  confReg_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  confReg_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  confReg_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  confReg_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  confReg_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  confReg_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  confReg_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  confReg_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  confReg_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  confReg_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  confReg_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  confReg_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  confReg_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  confReg_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  confReg_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  confReg_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  confReg_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  confReg_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  confReg_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  confReg_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  confReg_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  confReg_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  confReg_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  confReg_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  confReg_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  confReg_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  confReg_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  confReg_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  confReg_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  confReg_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  confReg_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  confReg_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  confReg_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  confReg_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  confReg_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  confReg_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  confReg_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  confReg_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  confReg_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  confReg_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  confReg_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  confReg_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  confReg_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  confReg_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  confReg_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  confReg_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  confReg_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  confReg_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  confReg_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  confReg_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  confReg_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  confReg_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  confReg_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  confReg_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  confReg_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  confReg_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  confReg_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  confReg_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  confReg_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  confReg_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  confReg_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  confReg_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  confReg_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  confReg_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  confReg_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  confReg_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  confReg_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  confReg_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  confReg_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  confReg_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  confReg_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  confReg_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  confReg_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  confReg_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  confReg_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  confReg_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  confReg_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  confReg_257 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  confReg_258 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  confReg_259 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  confReg_260 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  confReg_261 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  confReg_262 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  confReg_263 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  confReg_264 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  confReg_265 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  confReg_266 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  confReg_267 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  confReg_268 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  confReg_269 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  confReg_270 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  confReg_271 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  confReg_272 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  confReg_273 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  confReg_274 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  confReg_275 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  confReg_276 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  confReg_277 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  confReg_278 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  confReg_279 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  confReg_280 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  confReg_281 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  confReg_282 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  confReg_283 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  confReg_284 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  confReg_285 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  confReg_286 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  confReg_287 = _RAND_287[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MuxNInput_O0_C2_SCAOptSB(
  input  [1:0] io_in,
  input  [1:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [1:0] OPinMux_in; // @[MuxListTest.scala 108:26]
  wire  OPinMux_sel; // @[MuxListTest.scala 108:26]
  wire  OPinMux_o; // @[MuxListTest.scala 108:26]
  wire [1:0] chanMux_in; // @[MuxListTest.scala 129:26]
  wire  chanMux_sel; // @[MuxListTest.scala 129:26]
  wire  chanMux_o; // @[MuxListTest.scala 129:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire  _OPinMux_sel_T = io_config[0]; // @[MuxListTest.scala 121:33]
  wire  _chanMux_sel_T = io_config[0]; // @[MuxListTest.scala 143:33]
  wire [1:0] _chanMux_in_T = io_in; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[1]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[1] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux2C OPinMux ( // @[MuxListTest.scala 108:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux2C chanMux ( // @[MuxListTest.scala 129:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = 2'h0; // @[MuxListTest.scala 125:22]
  assign OPinMux_sel = io_config[0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = io_in; // @[MuxListTest.scala 145:30]
  assign chanMux_sel = io_config[0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[1] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O0_C3_SCAOptSB(
  input  [2:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire [1:0] _OPinMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 121:33]
  wire [1:0] _chanMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 143:33]
  wire [2:0] _chanMux_in_T = io_in; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[2]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = 4'h0; // @[MuxListTest.scala 125:22]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{1'd0}, io_in}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O0_C5_SCAOptSB(
  input  [4:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire [2:0] _OPinMux_sel_T = io_config[2:0]; // @[MuxListTest.scala 121:33]
  wire [2:0] _chanMux_sel_T = io_config[2:0]; // @[MuxListTest.scala 143:33]
  wire [4:0] _chanMux_in_T = io_in; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[3]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[3] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = 8'h0; // @[MuxListTest.scala 125:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O0_C4_SCAOptSB(
  input  [3:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire [1:0] _OPinMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 121:33]
  wire [1:0] _chanMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 143:33]
  wire [3:0] _chanMux_in_T = io_in; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[2]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = 4'h0; // @[MuxListTest.scala 125:22]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = io_in; // @[MuxListTest.scala 145:30]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O2_C3_SCAOptSB(
  input  [4:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire [1:0] _OPinMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 121:33]
  wire [1:0] _OPinMux_in_T = io_in[1:0]; // @[MuxListTest.scala 123:30]
  wire [1:0] _chanMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 143:33]
  wire [2:0] _chanMux_in_T = io_in[4:2]; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[2]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{2'd0}, io_in[1:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{1'd0}, io_in[4:2]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O2_C4_SCAOptSB(
  input  [5:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire [1:0] _OPinMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 121:33]
  wire [1:0] _OPinMux_in_T = io_in[1:0]; // @[MuxListTest.scala 123:30]
  wire [1:0] _chanMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 143:33]
  wire [3:0] _chanMux_in_T = io_in[5:2]; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[2]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{2'd0}, io_in[1:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = io_in[5:2]; // @[MuxListTest.scala 145:30]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O2_C2_SCAOptSB(
  input  [3:0] io_in,
  input  [1:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [1:0] OPinMux_in; // @[MuxListTest.scala 108:26]
  wire  OPinMux_sel; // @[MuxListTest.scala 108:26]
  wire  OPinMux_o; // @[MuxListTest.scala 108:26]
  wire [1:0] chanMux_in; // @[MuxListTest.scala 129:26]
  wire  chanMux_sel; // @[MuxListTest.scala 129:26]
  wire  chanMux_o; // @[MuxListTest.scala 129:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire  _OPinMux_sel_T = io_config[0]; // @[MuxListTest.scala 121:33]
  wire [1:0] _OPinMux_in_T = io_in[1:0]; // @[MuxListTest.scala 123:30]
  wire  _chanMux_sel_T = io_config[0]; // @[MuxListTest.scala 143:33]
  wire [1:0] _chanMux_in_T = io_in[3:2]; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[1]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[1] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux2C OPinMux ( // @[MuxListTest.scala 108:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux2C chanMux ( // @[MuxListTest.scala 129:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = io_in[1:0]; // @[MuxListTest.scala 123:30]
  assign OPinMux_sel = io_config[0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = io_in[3:2]; // @[MuxListTest.scala 145:30]
  assign chanMux_sel = io_config[0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[1] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O1_C3_SCAOptSB(
  input  [3:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire [1:0] _OPinMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 121:33]
  wire  _OPinMux_in_T = io_in[0]; // @[MuxListTest.scala 123:30]
  wire [1:0] _chanMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 143:33]
  wire [2:0] _chanMux_in_T = io_in[3:1]; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[2]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{3'd0}, io_in[0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{1'd0}, io_in[3:1]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O1_C2_SCAOptSB(
  input  [2:0] io_in,
  input  [1:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [1:0] OPinMux_in; // @[MuxListTest.scala 108:26]
  wire  OPinMux_sel; // @[MuxListTest.scala 108:26]
  wire  OPinMux_o; // @[MuxListTest.scala 108:26]
  wire [1:0] chanMux_in; // @[MuxListTest.scala 129:26]
  wire  chanMux_sel; // @[MuxListTest.scala 129:26]
  wire  chanMux_o; // @[MuxListTest.scala 129:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire  _OPinMux_sel_T = io_config[0]; // @[MuxListTest.scala 121:33]
  wire  _OPinMux_in_T = io_in[0]; // @[MuxListTest.scala 123:30]
  wire  _chanMux_sel_T = io_config[0]; // @[MuxListTest.scala 143:33]
  wire [1:0] _chanMux_in_T = io_in[2:1]; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[1]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[1] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux2C OPinMux ( // @[MuxListTest.scala 108:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux2C chanMux ( // @[MuxListTest.scala 129:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{1'd0}, io_in[0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = io_in[2:1]; // @[MuxListTest.scala 145:30]
  assign chanMux_sel = io_config[0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[1] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O4_C2_SCAOptSB(
  input  [5:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire [1:0] _OPinMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 121:33]
  wire [3:0] _OPinMux_in_T = io_in[3:0]; // @[MuxListTest.scala 123:30]
  wire [1:0] _chanMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 143:33]
  wire [1:0] _chanMux_in_T = io_in[5:4]; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[2]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = io_in[3:0]; // @[MuxListTest.scala 123:30]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in[5:4]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O3_C2_SCAOptSB(
  input  [4:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  wire [1:0] _OPinMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 121:33]
  wire [2:0] _OPinMux_in_T = io_in[2:0]; // @[MuxListTest.scala 123:30]
  wire [1:0] _chanMux_sel_T = io_config[1:0]; // @[MuxListTest.scala 143:33]
  wire [1:0] _chanMux_in_T = io_in[4:3]; // @[MuxListTest.scala 145:30]
  wire  _lbSBFlop_io_d_T = chanMux_o & OPinMux_o; // @[MuxListTest.scala 153:34]
  wire  _lbSBFlop_io_d_T_1 = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  wire  _lbCBMux_io_sa_T = io_config[2]; // @[MuxListTest.scala 157:28]
  wire  _lbCBMux_io_sa_T_1 = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  wire  _io_out_T = lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:39]
  wire  _io_out_T_1 = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{1'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in[4:3]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module Tile_11_0_EMPTY(
  input          clock,
  input          reset,
  input          IN_OPIN_N21936_32,
  input          IN_OPIN_N21937_33,
  input          IN_OPIN_N21938_34,
  input          IN_OPIN_N21939_35,
  input          IN_OPIN_N21940_36,
  input          IN_OPIN_N21941_37,
  input          IN_OPIN_N21942_38,
  input          IN_OPIN_N21943_39,
  input          IN_OPIN_N21944_40,
  input          IN_OPIN_N21945_41,
  input          IN_OPIN_N21946_42,
  input          IN_OPIN_N21947_43,
  input          IN_OPIN_N21948_44,
  input          IN_OPIN_N21949_45,
  input          IN_OPIN_N21950_46,
  input          IN_OPIN_N21951_47,
  input          IN_OPIN_N21952_48,
  input          IN_OPIN_N21953_49,
  input          IN_OPIN_N21954_50,
  input          IN_OPIN_N21955_51,
  input          IN_OPIN_N21956_52,
  input          IN_OPIN_N21957_53,
  input          IN_OPIN_N21958_54,
  input          IN_OPIN_N21959_55,
  input          IN_OPIN_N21960_56,
  input          IN_OPIN_N21961_57,
  input          IN_OPIN_N21962_58,
  input          IN_OPIN_N21963_59,
  input          IN_OPIN_N21964_60,
  input          IN_OPIN_N21965_61,
  input          IN_OPIN_N21966_62,
  input          IN_OPIN_N21967_63,
  input          IN_CHANX_N23428_6,
  input          IN_CHANX_N23430_14,
  input          IN_CHANX_N23432_22,
  input          IN_CHANX_N23434_30,
  input          IN_CHANX_N23436_38,
  input          IN_CHANX_N23438_46,
  input          IN_CHANX_N23440_54,
  input          IN_CHANX_N23442_62,
  input          IN_CHANX_N23444_70,
  input          IN_CHANX_N23446_78,
  input          IN_CHANX_N23462_0,
  input          IN_CHANX_N23464_8,
  input          IN_CHANX_N23466_16,
  input          IN_CHANX_N23468_24,
  input          IN_CHANX_N23470_32,
  input          IN_CHANX_N23472_40,
  input          IN_CHANX_N23474_48,
  input          IN_CHANX_N23476_56,
  input          IN_CHANX_N23478_64,
  input          IN_CHANX_N23480_72,
  input          IN_CHANX_N23482_80,
  input          IN_CHANX_N23496_2,
  input          IN_CHANX_N23498_10,
  input          IN_CHANX_N23500_18,
  input          IN_CHANX_N23502_26,
  input          IN_CHANX_N23504_34,
  input          IN_CHANX_N23506_42,
  input          IN_CHANX_N23508_50,
  input          IN_CHANX_N23510_58,
  input          IN_CHANX_N23512_66,
  input          IN_CHANX_N23514_74,
  input          IN_CHANX_N23516_82,
  input          IN_CHANX_N23518_86,
  input          IN_CHANX_N23520_90,
  input          IN_CHANX_N23522_94,
  input          IN_CHANX_N23524_98,
  input          IN_CHANX_N23526_102,
  input          IN_CHANX_N23528_106,
  input          IN_CHANX_N23530_4,
  input          IN_CHANX_N23532_12,
  input          IN_CHANX_N23534_20,
  input          IN_CHANX_N23536_28,
  input          IN_CHANX_N23538_36,
  input          IN_CHANX_N23540_44,
  input          IN_CHANX_N23542_52,
  input          IN_CHANX_N23544_60,
  input          IN_CHANX_N23546_68,
  input          IN_CHANX_N23548_76,
  input          IN_CHANX_N23550_84,
  input          IN_CHANX_N23552_88,
  input          IN_CHANX_N23554_92,
  input          IN_CHANX_N23556_96,
  input          IN_CHANX_N23558_100,
  input          IN_CHANX_N23560_104,
  input          IN_CHANY_N32497_1,
  input          IN_CHANY_N32499_3,
  input          IN_CHANY_N32501_5,
  input          IN_CHANY_N32503_7,
  input          IN_CHANY_N32505_9,
  input          IN_CHANY_N32507_11,
  input          IN_CHANY_N32509_13,
  input          IN_CHANY_N32511_15,
  input          IN_CHANY_N32513_17,
  input          IN_CHANY_N32515_19,
  input          IN_CHANY_N32517_21,
  input          IN_CHANY_N32519_23,
  input          IN_CHANY_N32521_25,
  input          IN_CHANY_N32523_27,
  input          IN_CHANY_N32525_29,
  input          IN_CHANY_N32527_31,
  input          IN_CHANY_N32529_33,
  input          IN_CHANY_N32531_35,
  input          IN_CHANY_N32533_37,
  input          IN_CHANY_N32535_39,
  input          IN_CHANY_N32537_41,
  input          IN_CHANY_N32539_43,
  input          IN_CHANY_N32541_45,
  input          IN_CHANY_N32543_47,
  input          IN_CHANY_N32545_49,
  input          IN_CHANY_N32547_51,
  input          IN_CHANY_N32549_53,
  input          IN_CHANY_N32551_55,
  input          IN_CHANY_N32553_57,
  input          IN_CHANY_N32555_59,
  input          IN_CHANY_N32557_61,
  input          IN_CHANY_N32559_63,
  input          IN_CHANY_N32561_65,
  input          IN_CHANY_N32563_67,
  input          IN_CHANY_N32565_69,
  input          IN_CHANY_N32567_71,
  input          IN_CHANY_N32569_73,
  input          IN_CHANY_N32571_75,
  input          IN_CHANY_N32573_77,
  input          IN_CHANY_N32575_79,
  input          IN_CHANY_N32577_81,
  input          IN_CHANY_N32579_83,
  input          IN_CHANY_N32581_85,
  input          IN_CHANY_N32583_87,
  input          IN_CHANY_N32585_89,
  input          IN_CHANY_N32587_91,
  input          IN_CHANY_N32589_93,
  input          IN_CHANY_N32591_95,
  input          IN_CHANY_N32593_97,
  input          IN_CHANY_N32595_99,
  input          IN_CHANY_N32597_101,
  input          IN_CHANY_N32599_103,
  input          IN_CHANY_N32601_105,
  input          IN_CHANY_N32603_107,
  output         OUT_CHANY_N32528_32,
  output         OUT_CHANY_N32584_88,
  output         OUT_CHANY_N32566_70,
  output         OUT_CHANX_N23429_7,
  output         OUT_CHANX_N23537_29,
  output         OUT_CHANX_N23553_89,
  output         OUT_CHANY_N32568_72,
  output         OUT_CHANX_N23523_95,
  output         OUT_CHANY_N32534_38,
  output         OUT_CHANY_N32586_90,
  output         OUT_CHANY_N32546_50,
  output         OUT_CHANY_N32512_16,
  output         OUT_CHANY_N32554_58,
  output         OUT_CHANX_N23505_35,
  output         OUT_CHANY_N32548_52,
  output         OUT_CHANX_N23543_53,
  output         OUT_CHANY_N32596_100,
  output         OUT_CHANY_N32594_98,
  output         OUT_CHANY_N32560_64,
  output         OUT_CHANX_N23521_91,
  output         OUT_CHANY_N32582_86,
  output         OUT_CHANY_N32598_102,
  output         OUT_CHANX_N23527_103,
  output         OUT_CHANX_N23551_85,
  output         OUT_CHANY_N32508_12,
  output         OUT_CHANY_N32570_74,
  output         OUT_CHANX_N23499_11,
  output         OUT_CHANY_N32502_6,
  output         OUT_CHANX_N23535_21,
  output         OUT_CHANX_N23525_99,
  output         OUT_CHANX_N23501_19,
  output         OUT_CHANY_N32580_84,
  output         OUT_CHANX_N23517_83,
  output         OUT_CHANX_N23531_5,
  output         OUT_CHANY_N32524_28,
  output         OUT_CHANY_N32532_36,
  output         OUT_CHANY_N32602_106,
  output         OUT_CHANX_N23477_57,
  output         OUT_CHANX_N23473_41,
  output         OUT_CHANX_N23479_65,
  output         OUT_CHANY_N32552_56,
  output         OUT_CHANX_N23555_93,
  output         OUT_CHANX_N23447_79,
  output         OUT_CHANY_N32592_96,
  output         OUT_CHANX_N23561_105,
  output         OUT_CHANY_N32522_26,
  output         OUT_CHANX_N23513_67,
  output         OUT_CHANY_N32510_14,
  output         OUT_CHANY_N32544_48,
  output         OUT_CHANX_N23431_15,
  output         OUT_CHANX_N23435_31,
  output         OUT_CHANX_N23503_27,
  output         OUT_CHANY_N32518_22,
  output         OUT_CHANX_N23463_1,
  output         OUT_CHANX_N23437_39,
  output         OUT_CHANY_N32530_34,
  output         OUT_CHANY_N32496_0,
  output         OUT_CHANX_N23529_107,
  output         OUT_CHANX_N23469_25,
  output         OUT_CHANY_N32588_92,
  output         OUT_CHANY_N32536_40,
  output         OUT_CHANY_N32574_78,
  output         OUT_CHANY_N32578_82,
  output         OUT_CHANX_N23475_49,
  output         OUT_CHANY_N32550_54,
  output         OUT_CHANX_N23443_63,
  output         OUT_CHANY_N32564_68,
  output         OUT_CHANX_N23467_17,
  output         OUT_CHANX_N23471_33,
  output         OUT_CHANX_N23433_23,
  output         OUT_CHANY_N32558_62,
  output         OUT_CHANX_N23559_101,
  output         OUT_CHANY_N32516_20,
  output         OUT_CHANX_N23549_77,
  output         OUT_CHANY_N32526_30,
  output         OUT_CHANY_N32500_4,
  output         OUT_CHANX_N23445_71,
  output         OUT_CHANY_N32498_2,
  output         OUT_CHANX_N23481_73,
  output         OUT_CHANY_N32540_44,
  output         OUT_CHANX_N23539_37,
  output         OUT_CHANY_N32506_10,
  output         OUT_CHANX_N23465_9,
  output         OUT_CHANX_N23483_81,
  output         OUT_CHANX_N23439_47,
  output         OUT_CHANY_N32576_80,
  output         OUT_CHANX_N23545_61,
  output         OUT_CHANX_N23515_75,
  output         OUT_CHANY_N32520_24,
  output         OUT_CHANX_N23497_3,
  output         OUT_CHANX_N23509_51,
  output         OUT_CHANX_N23541_45,
  output         OUT_CHANY_N32538_42,
  output         OUT_CHANY_N32542_46,
  output         OUT_CHANY_N32572_76,
  output         OUT_CHANX_N23507_43,
  output         OUT_CHANY_N32504_8,
  output         OUT_CHANY_N32600_104,
  output         OUT_CHANY_N32556_60,
  output         OUT_CHANY_N32590_94,
  output         OUT_CHANY_N32514_18,
  output         OUT_CHANY_N32562_66,
  output         OUT_CHANX_N23511_59,
  output         OUT_CHANX_N23441_55,
  output         OUT_CHANX_N23519_87,
  output         OUT_CHANX_N23533_13,
  output         OUT_CHANX_N23557_97,
  output         OUT_CHANX_N23547_69,
  output [282:0] ioConf_confOut,
  input  [15:0]  ioConf_scan_in,
  input          ioConf_scan_en,
  output [15:0]  ioConf_scan_out,
  input          ioConf_scan_ioLatchEnb,
  input          ctrlSignals_gndBlkOuts,
  input          ctrlSignals_loopBreak,
  input          ctrlSignals_arst,
  input          ctrlSignals_confClock,
  input          ctrlSignals_constClock
);
  wire  configBlock_clock; // @[TileFull.scala 67:31]
  wire  configBlock_reset; // @[TileFull.scala 67:31]
  wire [287:0] configBlock_ioBundle_confOut; // @[TileFull.scala 67:31]
  wire [15:0] configBlock_ioBundle_scan_in; // @[TileFull.scala 67:31]
  wire  configBlock_ioBundle_scan_en; // @[TileFull.scala 67:31]
  wire [15:0] configBlock_ioBundle_scan_out; // @[TileFull.scala 67:31]
  wire  configBlock_ioBundle_scan_ioLatchEnb; // @[TileFull.scala 67:31]
  wire [1:0] SBMux_C7_N23429_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C7_N23429_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C7_N23429_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C7_N23429_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C7_N23429_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C7_N23429_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C7_N23429_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C15_N23431_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C15_N23431_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C15_N23431_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C15_N23431_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C15_N23431_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C15_N23431_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C15_N23431_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C23_N23433_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C23_N23433_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C23_N23433_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C23_N23433_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C23_N23433_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C23_N23433_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C23_N23433_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C31_N23435_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C31_N23435_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C31_N23435_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C31_N23435_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C31_N23435_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C31_N23435_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C31_N23435_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C39_N23437_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C39_N23437_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C39_N23437_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C39_N23437_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C39_N23437_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C39_N23437_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C39_N23437_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C47_N23439_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C47_N23439_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C47_N23439_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C47_N23439_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C47_N23439_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C47_N23439_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C47_N23439_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C55_N23441_O_0_C_5_io_in; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C55_N23441_O_0_C_5_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C55_N23441_O_0_C_5_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C55_N23441_O_0_C_5_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C55_N23441_O_0_C_5_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C55_N23441_O_0_C_5_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C55_N23441_O_0_C_5_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C63_N23443_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C63_N23443_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C63_N23443_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C63_N23443_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C63_N23443_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C63_N23443_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C63_N23443_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C71_N23445_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C71_N23445_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C71_N23445_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C71_N23445_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C71_N23445_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C71_N23445_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C71_N23445_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C79_N23447_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C79_N23447_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C79_N23447_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C79_N23447_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C79_N23447_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C79_N23447_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C79_N23447_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C1_N23463_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C1_N23463_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C1_N23463_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C1_N23463_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C1_N23463_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C1_N23463_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C1_N23463_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C9_N23465_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C9_N23465_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C9_N23465_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C9_N23465_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C9_N23465_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C9_N23465_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C9_N23465_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C17_N23467_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C17_N23467_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C17_N23467_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C17_N23467_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C17_N23467_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C17_N23467_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C17_N23467_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C25_N23469_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C25_N23469_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C25_N23469_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C25_N23469_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C25_N23469_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C25_N23469_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C25_N23469_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C33_N23471_O_0_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C33_N23471_O_0_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C33_N23471_O_0_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C33_N23471_O_0_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C33_N23471_O_0_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C33_N23471_O_0_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C33_N23471_O_0_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C41_N23473_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C41_N23473_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C41_N23473_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C41_N23473_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C41_N23473_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C41_N23473_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C41_N23473_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C49_N23475_O_0_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C49_N23475_O_0_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C49_N23475_O_0_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C49_N23475_O_0_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C49_N23475_O_0_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C49_N23475_O_0_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C49_N23475_O_0_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C57_N23477_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C57_N23477_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C57_N23477_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C57_N23477_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C57_N23477_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C57_N23477_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C57_N23477_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C65_N23479_O_0_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C65_N23479_O_0_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C65_N23479_O_0_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C65_N23479_O_0_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C65_N23479_O_0_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C65_N23479_O_0_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C65_N23479_O_0_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C73_N23481_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C73_N23481_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C73_N23481_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C73_N23481_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C73_N23481_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C73_N23481_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C73_N23481_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C81_N23483_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C81_N23483_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C81_N23483_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C81_N23483_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C81_N23483_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C81_N23483_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C81_N23483_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C3_N23497_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C3_N23497_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C3_N23497_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C3_N23497_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C3_N23497_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C3_N23497_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C3_N23497_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C11_N23499_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C11_N23499_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C11_N23499_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C11_N23499_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C11_N23499_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C11_N23499_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C11_N23499_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C19_N23501_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C19_N23501_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C19_N23501_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C19_N23501_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C19_N23501_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C19_N23501_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C19_N23501_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C27_N23503_O_0_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C27_N23503_O_0_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C27_N23503_O_0_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C27_N23503_O_0_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C27_N23503_O_0_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C27_N23503_O_0_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C27_N23503_O_0_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C35_N23505_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C35_N23505_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C35_N23505_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C35_N23505_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C35_N23505_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C35_N23505_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C35_N23505_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C43_N23507_O_0_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C43_N23507_O_0_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C43_N23507_O_0_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C43_N23507_O_0_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C43_N23507_O_0_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C43_N23507_O_0_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C43_N23507_O_0_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C51_N23509_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C51_N23509_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C51_N23509_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C51_N23509_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C51_N23509_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C51_N23509_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C51_N23509_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C59_N23511_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C59_N23511_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C59_N23511_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C59_N23511_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C59_N23511_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C59_N23511_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C59_N23511_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C67_N23513_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C67_N23513_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C67_N23513_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C67_N23513_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C67_N23513_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C67_N23513_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C67_N23513_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C75_N23515_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C75_N23515_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C75_N23515_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C75_N23515_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C75_N23515_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C75_N23515_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C75_N23515_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C83_N23517_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C83_N23517_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C83_N23517_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C83_N23517_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C83_N23517_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C83_N23517_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C83_N23517_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C87_N23519_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C87_N23519_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C87_N23519_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C87_N23519_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C87_N23519_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C87_N23519_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C87_N23519_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C91_N23521_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C91_N23521_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C91_N23521_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C91_N23521_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C91_N23521_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C91_N23521_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C91_N23521_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C95_N23523_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C95_N23523_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C95_N23523_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C95_N23523_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C95_N23523_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C95_N23523_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C95_N23523_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C99_N23525_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C99_N23525_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C99_N23525_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C99_N23525_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C99_N23525_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C99_N23525_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C99_N23525_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C103_N23527_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C103_N23527_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C103_N23527_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C103_N23527_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C103_N23527_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C103_N23527_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C103_N23527_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C107_N23529_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C107_N23529_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C107_N23529_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C107_N23529_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C107_N23529_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C107_N23529_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C107_N23529_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C5_N23531_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C5_N23531_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C5_N23531_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C5_N23531_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C5_N23531_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C5_N23531_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C5_N23531_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C13_N23533_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C13_N23533_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C13_N23533_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C13_N23533_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C13_N23533_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C13_N23533_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C13_N23533_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C21_N23535_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C21_N23535_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C21_N23535_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C21_N23535_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C21_N23535_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C21_N23535_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C21_N23535_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C29_N23537_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C29_N23537_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C29_N23537_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C29_N23537_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C29_N23537_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C29_N23537_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C29_N23537_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C37_N23539_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C37_N23539_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C37_N23539_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C37_N23539_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C37_N23539_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C37_N23539_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C37_N23539_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C45_N23541_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C45_N23541_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C45_N23541_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C45_N23541_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C45_N23541_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C45_N23541_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C45_N23541_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C53_N23543_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C53_N23543_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C53_N23543_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C53_N23543_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C53_N23543_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C53_N23543_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C53_N23543_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C61_N23545_O_0_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C61_N23545_O_0_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C61_N23545_O_0_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C61_N23545_O_0_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C61_N23545_O_0_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C61_N23545_O_0_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C61_N23545_O_0_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C69_N23547_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C69_N23547_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C69_N23547_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C69_N23547_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C69_N23547_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C69_N23547_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C69_N23547_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C77_N23549_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C77_N23549_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C77_N23549_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C77_N23549_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C77_N23549_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C77_N23549_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C77_N23549_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C85_N23551_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C85_N23551_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C85_N23551_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C85_N23551_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C85_N23551_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C85_N23551_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C85_N23551_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C89_N23553_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C89_N23553_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C89_N23553_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C89_N23553_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C89_N23553_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C89_N23553_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C89_N23553_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C93_N23555_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C93_N23555_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C93_N23555_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C93_N23555_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C93_N23555_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C93_N23555_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C93_N23555_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C97_N23557_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C97_N23557_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C97_N23557_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C97_N23557_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C97_N23557_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C97_N23557_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C97_N23557_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C101_N23559_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C101_N23559_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C101_N23559_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C101_N23559_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C101_N23559_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C101_N23559_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C101_N23559_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C105_N23561_O_0_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C105_N23561_O_0_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C105_N23561_O_0_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C105_N23561_O_0_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C105_N23561_O_0_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C105_N23561_O_0_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C105_N23561_O_0_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C0_N32496_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C0_N32496_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C0_N32496_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C0_N32496_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C0_N32496_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C0_N32496_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C0_N32496_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C2_N32498_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C2_N32498_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C2_N32498_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C2_N32498_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C2_N32498_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C2_N32498_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C2_N32498_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C4_N32500_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C4_N32500_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C4_N32500_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C4_N32500_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C4_N32500_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C4_N32500_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C4_N32500_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C6_N32502_O_2_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C6_N32502_O_2_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C6_N32502_O_2_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C6_N32502_O_2_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C6_N32502_O_2_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C6_N32502_O_2_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C6_N32502_O_2_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C8_N32504_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C8_N32504_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C8_N32504_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C8_N32504_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C8_N32504_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C8_N32504_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C8_N32504_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C10_N32506_O_2_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C10_N32506_O_2_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C10_N32506_O_2_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C10_N32506_O_2_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C10_N32506_O_2_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C10_N32506_O_2_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C10_N32506_O_2_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C12_N32508_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C12_N32508_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C12_N32508_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C12_N32508_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C12_N32508_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C12_N32508_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C12_N32508_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C14_N32510_O_2_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C14_N32510_O_2_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C14_N32510_O_2_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C14_N32510_O_2_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C14_N32510_O_2_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C14_N32510_O_2_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C14_N32510_O_2_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C16_N32512_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C16_N32512_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C16_N32512_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C16_N32512_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C16_N32512_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C16_N32512_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C16_N32512_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C18_N32514_O_2_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C18_N32514_O_2_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C18_N32514_O_2_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C18_N32514_O_2_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C18_N32514_O_2_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C18_N32514_O_2_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C18_N32514_O_2_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C20_N32516_O_2_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C20_N32516_O_2_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C20_N32516_O_2_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C20_N32516_O_2_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C20_N32516_O_2_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C20_N32516_O_2_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C20_N32516_O_2_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C22_N32518_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C22_N32518_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C22_N32518_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C22_N32518_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C22_N32518_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C22_N32518_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C22_N32518_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C24_N32520_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C24_N32520_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C24_N32520_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C24_N32520_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C24_N32520_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C24_N32520_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C24_N32520_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C26_N32522_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C26_N32522_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C26_N32522_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C26_N32522_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C26_N32522_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C26_N32522_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C26_N32522_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C28_N32524_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C28_N32524_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C28_N32524_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C28_N32524_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C28_N32524_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C28_N32524_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C28_N32524_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C30_N32526_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C30_N32526_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C30_N32526_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C30_N32526_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C30_N32526_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C30_N32526_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C30_N32526_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C32_N32528_O_2_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C32_N32528_O_2_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C32_N32528_O_2_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C32_N32528_O_2_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C32_N32528_O_2_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C32_N32528_O_2_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C32_N32528_O_2_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C34_N32530_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C34_N32530_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C34_N32530_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C34_N32530_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C34_N32530_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C34_N32530_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C34_N32530_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C36_N32532_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C36_N32532_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C36_N32532_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C36_N32532_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C36_N32532_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C36_N32532_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C36_N32532_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C38_N32534_O_2_C_4_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C38_N32534_O_2_C_4_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C38_N32534_O_2_C_4_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C38_N32534_O_2_C_4_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C38_N32534_O_2_C_4_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C38_N32534_O_2_C_4_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C38_N32534_O_2_C_4_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C40_N32536_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C40_N32536_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C40_N32536_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C40_N32536_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C40_N32536_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C40_N32536_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C40_N32536_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C42_N32538_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C42_N32538_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C42_N32538_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C42_N32538_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C42_N32538_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C42_N32538_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C42_N32538_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C44_N32540_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C44_N32540_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C44_N32540_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C44_N32540_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C44_N32540_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C44_N32540_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C44_N32540_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C46_N32542_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C46_N32542_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C46_N32542_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C46_N32542_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C46_N32542_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C46_N32542_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C46_N32542_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C48_N32544_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C48_N32544_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C48_N32544_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C48_N32544_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C48_N32544_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C48_N32544_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C48_N32544_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C50_N32546_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C50_N32546_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C50_N32546_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C50_N32546_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C50_N32546_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C50_N32546_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C50_N32546_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C52_N32548_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C52_N32548_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C52_N32548_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C52_N32548_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C52_N32548_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C52_N32548_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C52_N32548_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C54_N32550_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C54_N32550_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C54_N32550_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C54_N32550_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C54_N32550_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C54_N32550_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C54_N32550_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C56_N32552_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C56_N32552_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C56_N32552_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C56_N32552_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C56_N32552_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C56_N32552_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C56_N32552_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C58_N32554_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C58_N32554_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C58_N32554_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C58_N32554_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C58_N32554_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C58_N32554_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C58_N32554_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C60_N32556_O_2_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C60_N32556_O_2_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C60_N32556_O_2_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C60_N32556_O_2_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C60_N32556_O_2_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C60_N32556_O_2_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C60_N32556_O_2_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C62_N32558_O_1_C_3_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C62_N32558_O_1_C_3_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C62_N32558_O_1_C_3_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C62_N32558_O_1_C_3_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C62_N32558_O_1_C_3_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C62_N32558_O_1_C_3_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C62_N32558_O_1_C_3_io_arst; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C64_N32560_O_1_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C64_N32560_O_1_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C64_N32560_O_1_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C64_N32560_O_1_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C64_N32560_O_1_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C64_N32560_O_1_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C64_N32560_O_1_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C66_N32562_O_4_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C66_N32562_O_4_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C66_N32562_O_4_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C66_N32562_O_4_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C66_N32562_O_4_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C66_N32562_O_4_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C66_N32562_O_4_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C68_N32564_O_4_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C68_N32564_O_4_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C68_N32564_O_4_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C68_N32564_O_4_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C68_N32564_O_4_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C68_N32564_O_4_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C68_N32564_O_4_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C70_N32566_O_4_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C70_N32566_O_4_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C70_N32566_O_4_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C70_N32566_O_4_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C70_N32566_O_4_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C70_N32566_O_4_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C70_N32566_O_4_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C72_N32568_O_4_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C72_N32568_O_4_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C72_N32568_O_4_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C72_N32568_O_4_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C72_N32568_O_4_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C72_N32568_O_4_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C72_N32568_O_4_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C74_N32570_O_4_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C74_N32570_O_4_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C74_N32570_O_4_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C74_N32570_O_4_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C74_N32570_O_4_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C74_N32570_O_4_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C74_N32570_O_4_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C76_N32572_O_4_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C76_N32572_O_4_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C76_N32572_O_4_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C76_N32572_O_4_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C76_N32572_O_4_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C76_N32572_O_4_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C76_N32572_O_4_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C78_N32574_O_4_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C78_N32574_O_4_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C78_N32574_O_4_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C78_N32574_O_4_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C78_N32574_O_4_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C78_N32574_O_4_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C78_N32574_O_4_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [5:0] SBMux_C80_N32576_O_4_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C80_N32576_O_4_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C80_N32576_O_4_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C80_N32576_O_4_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C80_N32576_O_4_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C80_N32576_O_4_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C80_N32576_O_4_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C82_N32578_O_3_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C82_N32578_O_3_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C82_N32578_O_3_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C82_N32578_O_3_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C82_N32578_O_3_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C82_N32578_O_3_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C82_N32578_O_3_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C84_N32580_O_3_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C84_N32580_O_3_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C84_N32580_O_3_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C84_N32580_O_3_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C84_N32580_O_3_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C84_N32580_O_3_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C84_N32580_O_3_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C86_N32582_O_3_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C86_N32582_O_3_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C86_N32582_O_3_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C86_N32582_O_3_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C86_N32582_O_3_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C86_N32582_O_3_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C86_N32582_O_3_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C88_N32584_O_3_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C88_N32584_O_3_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C88_N32584_O_3_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C88_N32584_O_3_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C88_N32584_O_3_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C88_N32584_O_3_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C88_N32584_O_3_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C90_N32586_O_3_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C90_N32586_O_3_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C90_N32586_O_3_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C90_N32586_O_3_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C90_N32586_O_3_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C90_N32586_O_3_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C90_N32586_O_3_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [4:0] SBMux_C92_N32588_O_3_C_2_io_in; // @[TileFull.scala 146:27]
  wire [2:0] SBMux_C92_N32588_O_3_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C92_N32588_O_3_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C92_N32588_O_3_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C92_N32588_O_3_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C92_N32588_O_3_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C92_N32588_O_3_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C94_N32590_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C94_N32590_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C94_N32590_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C94_N32590_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C94_N32590_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C94_N32590_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C94_N32590_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C96_N32592_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C96_N32592_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C96_N32592_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C96_N32592_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C96_N32592_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C96_N32592_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C96_N32592_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C98_N32594_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C98_N32594_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C98_N32594_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C98_N32594_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C98_N32594_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C98_N32594_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C98_N32594_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C100_N32596_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C100_N32596_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C100_N32596_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C100_N32596_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C100_N32596_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C100_N32596_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C100_N32596_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C102_N32598_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C102_N32598_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C102_N32598_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C102_N32598_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C102_N32598_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C102_N32598_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C102_N32598_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C104_N32600_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C104_N32600_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C104_N32600_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C104_N32600_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C104_N32600_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C104_N32600_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C104_N32600_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [3:0] SBMux_C106_N32602_O_2_C_2_io_in; // @[TileFull.scala 146:27]
  wire [1:0] SBMux_C106_N32602_O_2_C_2_io_config; // @[TileFull.scala 146:27]
  wire  SBMux_C106_N32602_O_2_C_2_io_out; // @[TileFull.scala 146:27]
  wire  SBMux_C106_N32602_O_2_C_2_io_loopBreak; // @[TileFull.scala 146:27]
  wire  SBMux_C106_N32602_O_2_C_2_io_ioGndBle; // @[TileFull.scala 146:27]
  wire  SBMux_C106_N32602_O_2_C_2_io_cnstClk; // @[TileFull.scala 146:27]
  wire  SBMux_C106_N32602_O_2_C_2_io_arst; // @[TileFull.scala 146:27]
  wire [1:0] _SBMux_C7_N23429_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[1:0]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C15_N23431_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[4:2]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C23_N23433_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[7:5]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C31_N23435_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[10:8]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C39_N23437_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[13:11]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C47_N23439_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[16:14]; // @[TileFull.scala 156:60]
  wire [3:0] _SBMux_C55_N23441_O_0_C_5_io_config_T = configBlock_ioBundle_confOut[20:17]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C63_N23443_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[23:21]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C71_N23445_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[25:24]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C79_N23447_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[27:26]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C1_N23463_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[29:28]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C9_N23465_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[32:30]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C17_N23467_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[35:33]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C25_N23469_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[38:36]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C33_N23471_O_0_C_4_io_config_T = configBlock_ioBundle_confOut[41:39]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C41_N23473_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[44:42]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C49_N23475_O_0_C_4_io_config_T = configBlock_ioBundle_confOut[47:45]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C57_N23477_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[50:48]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C65_N23479_O_0_C_4_io_config_T = configBlock_ioBundle_confOut[53:51]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C73_N23481_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[55:54]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C81_N23483_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[57:56]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C3_N23497_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[60:58]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C11_N23499_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[63:61]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C19_N23501_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[66:64]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C27_N23503_O_0_C_4_io_config_T = configBlock_ioBundle_confOut[69:67]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C35_N23505_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[72:70]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C43_N23507_O_0_C_4_io_config_T = configBlock_ioBundle_confOut[75:73]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C51_N23509_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[77:76]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C59_N23511_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[80:78]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C67_N23513_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[82:81]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C75_N23515_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[84:83]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C83_N23517_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[86:85]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C87_N23519_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[88:87]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C91_N23521_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[90:89]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C95_N23523_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[92:91]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C99_N23525_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[94:93]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C103_N23527_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[96:95]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C107_N23529_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[98:97]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C5_N23531_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[100:99]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C13_N23533_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[102:101]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C21_N23535_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[105:103]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C29_N23537_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[107:106]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C37_N23539_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[110:108]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C45_N23541_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[112:111]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C53_N23543_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[115:113]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C61_N23545_O_0_C_3_io_config_T = configBlock_ioBundle_confOut[118:116]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C69_N23547_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[120:119]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C77_N23549_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[122:121]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C85_N23551_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[124:123]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C89_N23553_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[126:125]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C93_N23555_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[128:127]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C97_N23557_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[130:129]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C101_N23559_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[132:131]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C105_N23561_O_0_C_2_io_config_T = configBlock_ioBundle_confOut[134:133]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C0_N32496_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[137:135]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C2_N32498_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[140:138]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C4_N32500_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[143:141]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C6_N32502_O_2_C_4_io_config_T = configBlock_ioBundle_confOut[146:144]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C8_N32504_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[149:147]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C10_N32506_O_2_C_4_io_config_T = configBlock_ioBundle_confOut[152:150]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C12_N32508_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[155:153]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C14_N32510_O_2_C_4_io_config_T = configBlock_ioBundle_confOut[158:156]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C16_N32512_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[161:159]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C18_N32514_O_2_C_4_io_config_T = configBlock_ioBundle_confOut[164:162]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C20_N32516_O_2_C_4_io_config_T = configBlock_ioBundle_confOut[167:165]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C22_N32518_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[170:168]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C24_N32520_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[172:171]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C26_N32522_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[175:173]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C28_N32524_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[177:176]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C30_N32526_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[179:178]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C32_N32528_O_2_C_4_io_config_T = configBlock_ioBundle_confOut[182:180]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C34_N32530_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[185:183]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C36_N32532_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[188:186]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C38_N32534_O_2_C_4_io_config_T = configBlock_ioBundle_confOut[191:189]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C40_N32536_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[193:192]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C42_N32538_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[196:194]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C44_N32540_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[199:197]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C46_N32542_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[202:200]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C48_N32544_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[205:203]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C50_N32546_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[208:206]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C52_N32548_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[211:209]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C54_N32550_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[213:212]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C56_N32552_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[216:214]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C58_N32554_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[218:217]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C60_N32556_O_2_C_3_io_config_T = configBlock_ioBundle_confOut[221:219]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C62_N32558_O_1_C_3_io_config_T = configBlock_ioBundle_confOut[224:222]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C64_N32560_O_1_C_2_io_config_T = configBlock_ioBundle_confOut[226:225]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C66_N32562_O_4_C_2_io_config_T = configBlock_ioBundle_confOut[229:227]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C68_N32564_O_4_C_2_io_config_T = configBlock_ioBundle_confOut[232:230]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C70_N32566_O_4_C_2_io_config_T = configBlock_ioBundle_confOut[235:233]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C72_N32568_O_4_C_2_io_config_T = configBlock_ioBundle_confOut[238:236]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C74_N32570_O_4_C_2_io_config_T = configBlock_ioBundle_confOut[241:239]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C76_N32572_O_4_C_2_io_config_T = configBlock_ioBundle_confOut[244:242]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C78_N32574_O_4_C_2_io_config_T = configBlock_ioBundle_confOut[247:245]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C80_N32576_O_4_C_2_io_config_T = configBlock_ioBundle_confOut[250:248]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C82_N32578_O_3_C_2_io_config_T = configBlock_ioBundle_confOut[253:251]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C84_N32580_O_3_C_2_io_config_T = configBlock_ioBundle_confOut[256:254]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C86_N32582_O_3_C_2_io_config_T = configBlock_ioBundle_confOut[259:257]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C88_N32584_O_3_C_2_io_config_T = configBlock_ioBundle_confOut[262:260]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C90_N32586_O_3_C_2_io_config_T = configBlock_ioBundle_confOut[265:263]; // @[TileFull.scala 156:60]
  wire [2:0] _SBMux_C92_N32588_O_3_C_2_io_config_T = configBlock_ioBundle_confOut[268:266]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C94_N32590_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[270:269]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C96_N32592_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[272:271]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C98_N32594_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[274:273]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C100_N32596_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[276:275]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C102_N32598_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[278:277]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C104_N32600_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[280:279]; // @[TileFull.scala 156:60]
  wire [1:0] _SBMux_C106_N32602_O_2_C_2_io_config_T = configBlock_ioBundle_confOut[282:281]; // @[TileFull.scala 156:60]
  wire  _SBMux_C7_N23429_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32569_73; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C7_N23429_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32529_33; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C7_N23429_O_0_C_2_io_in_T = {IN_CHANY_N32569_73,IN_CHANY_N32529_33}; // @[TileFull.scala 207:13]
  wire  _SBMux_C15_N23431_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32601_105; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C15_N23431_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32571_75; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C15_N23431_O_0_C_3_io_in_hi = {IN_CHANY_N32601_105,IN_CHANY_N32571_75}; // @[TileFull.scala 207:13]
  wire  _SBMux_C15_N23431_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32509_13; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C15_N23431_O_0_C_3_io_in_T = {IN_CHANY_N32601_105,IN_CHANY_N32571_75,IN_CHANY_N32509_13}; // @[TileFull.scala 207:13]
  wire  _SBMux_C23_N23433_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32581_85; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C23_N23433_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32575_79; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C23_N23433_O_0_C_3_io_in_hi = {IN_CHANY_N32581_85,IN_CHANY_N32575_79}; // @[TileFull.scala 207:13]
  wire  _SBMux_C23_N23433_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32505_9; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C23_N23433_O_0_C_3_io_in_T = {IN_CHANY_N32581_85,IN_CHANY_N32575_79,IN_CHANY_N32505_9}; // @[TileFull.scala 207:13]
  wire  _SBMux_C31_N23435_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32591_95; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C31_N23435_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32571_75; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C31_N23435_O_0_C_3_io_in_hi = {IN_CHANY_N32591_95,IN_CHANY_N32571_75}; // @[TileFull.scala 207:13]
  wire  _SBMux_C31_N23435_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32561_65; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C31_N23435_O_0_C_3_io_in_T = {IN_CHANY_N32591_95,IN_CHANY_N32571_75,IN_CHANY_N32561_65}; // @[TileFull.scala 207:13]
  wire  _SBMux_C39_N23437_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32583_87; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C39_N23437_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32563_67; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C39_N23437_O_0_C_3_io_in_hi = {IN_CHANY_N32583_87,IN_CHANY_N32563_67}; // @[TileFull.scala 207:13]
  wire  _SBMux_C39_N23437_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32513_17; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C39_N23437_O_0_C_3_io_in_T = {IN_CHANY_N32583_87,IN_CHANY_N32563_67,IN_CHANY_N32513_17}; // @[TileFull.scala 207:13]
  wire  _SBMux_C47_N23439_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32585_89; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C47_N23439_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32573_77; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C47_N23439_O_0_C_3_io_in_hi = {IN_CHANY_N32585_89,IN_CHANY_N32573_77}; // @[TileFull.scala 207:13]
  wire  _SBMux_C47_N23439_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32535_39; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C47_N23439_O_0_C_3_io_in_T = {IN_CHANY_N32585_89,IN_CHANY_N32573_77,IN_CHANY_N32535_39}; // @[TileFull.scala 207:13]
  wire  _SBMux_C55_N23441_O_0_C_5_io_in_WIRE_1 = IN_CHANY_N32567_71; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C55_N23441_O_0_C_5_io_in_WIRE_0 = IN_CHANY_N32533_37; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C55_N23441_O_0_C_5_io_in_lo = {IN_CHANY_N32567_71,IN_CHANY_N32533_37}; // @[TileFull.scala 207:13]
  wire  _SBMux_C55_N23441_O_0_C_5_io_in_WIRE_4 = IN_CHANY_N32599_103; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C55_N23441_O_0_C_5_io_in_WIRE_3 = IN_CHANY_N32583_87; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C55_N23441_O_0_C_5_io_in_hi_hi = {IN_CHANY_N32599_103,IN_CHANY_N32583_87}; // @[TileFull.scala 207:13]
  wire  _SBMux_C55_N23441_O_0_C_5_io_in_WIRE_2 = IN_CHANY_N32577_81; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C55_N23441_O_0_C_5_io_in_hi = {IN_CHANY_N32599_103,IN_CHANY_N32583_87,IN_CHANY_N32577_81}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C55_N23441_O_0_C_5_io_in_T = {IN_CHANY_N32599_103,IN_CHANY_N32583_87,IN_CHANY_N32577_81,
    IN_CHANY_N32567_71,IN_CHANY_N32533_37}; // @[TileFull.scala 207:13]
  wire  _SBMux_C63_N23443_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32603_107; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C63_N23443_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32563_67; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C63_N23443_O_0_C_3_io_in_hi = {IN_CHANY_N32603_107,IN_CHANY_N32563_67}; // @[TileFull.scala 207:13]
  wire  _SBMux_C63_N23443_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32511_15; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C63_N23443_O_0_C_3_io_in_T = {IN_CHANY_N32603_107,IN_CHANY_N32563_67,IN_CHANY_N32511_15}; // @[TileFull.scala 207:13]
  wire  _SBMux_C71_N23445_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32599_103; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C71_N23445_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32567_71; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C71_N23445_O_0_C_2_io_in_T = {IN_CHANY_N32599_103,IN_CHANY_N32567_71}; // @[TileFull.scala 207:13]
  wire  _SBMux_C79_N23447_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32597_101; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C79_N23447_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32563_67; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C79_N23447_O_0_C_2_io_in_T = {IN_CHANY_N32597_101,IN_CHANY_N32563_67}; // @[TileFull.scala 207:13]
  wire  _SBMux_C1_N23463_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32575_79; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C1_N23463_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32531_35; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C1_N23463_O_0_C_2_io_in_T = {IN_CHANY_N32575_79,IN_CHANY_N32531_35}; // @[TileFull.scala 207:13]
  wire  _SBMux_C9_N23465_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32591_95; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C9_N23465_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32577_81; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C9_N23465_O_0_C_3_io_in_hi = {IN_CHANY_N32591_95,IN_CHANY_N32577_81}; // @[TileFull.scala 207:13]
  wire  _SBMux_C9_N23465_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32501_5; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C9_N23465_O_0_C_3_io_in_T = {IN_CHANY_N32591_95,IN_CHANY_N32577_81,IN_CHANY_N32501_5}; // @[TileFull.scala 207:13]
  wire  _SBMux_C17_N23467_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32589_93; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C17_N23467_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32577_81; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C17_N23467_O_0_C_3_io_in_hi = {IN_CHANY_N32589_93,IN_CHANY_N32577_81}; // @[TileFull.scala 207:13]
  wire  _SBMux_C17_N23467_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32559_63; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C17_N23467_O_0_C_3_io_in_T = {IN_CHANY_N32589_93,IN_CHANY_N32577_81,IN_CHANY_N32559_63}; // @[TileFull.scala 207:13]
  wire  _SBMux_C25_N23469_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32597_101; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C25_N23469_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32565_69; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C25_N23469_O_0_C_3_io_in_hi = {IN_CHANY_N32597_101,IN_CHANY_N32565_69}; // @[TileFull.scala 207:13]
  wire  _SBMux_C25_N23469_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32555_59; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C25_N23469_O_0_C_3_io_in_T = {IN_CHANY_N32597_101,IN_CHANY_N32565_69,IN_CHANY_N32555_59}; // @[TileFull.scala 207:13]
  wire  _SBMux_C33_N23471_O_0_C_4_io_in_WIRE_1 = IN_CHANY_N32573_77; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C33_N23471_O_0_C_4_io_in_WIRE_0 = IN_CHANY_N32551_55; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C33_N23471_O_0_C_4_io_in_lo = {IN_CHANY_N32573_77,IN_CHANY_N32551_55}; // @[TileFull.scala 207:13]
  wire  _SBMux_C33_N23471_O_0_C_4_io_in_WIRE_3 = IN_CHANY_N32593_97; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C33_N23471_O_0_C_4_io_in_WIRE_2 = IN_CHANY_N32585_89; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C33_N23471_O_0_C_4_io_in_hi = {IN_CHANY_N32593_97,IN_CHANY_N32585_89}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C33_N23471_O_0_C_4_io_in_T = {IN_CHANY_N32593_97,IN_CHANY_N32585_89,IN_CHANY_N32573_77,
    IN_CHANY_N32551_55}; // @[TileFull.scala 207:13]
  wire  _SBMux_C41_N23473_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32581_85; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C41_N23473_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32565_69; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C41_N23473_O_0_C_3_io_in_hi = {IN_CHANY_N32581_85,IN_CHANY_N32565_69}; // @[TileFull.scala 207:13]
  wire  _SBMux_C41_N23473_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32541_45; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C41_N23473_O_0_C_3_io_in_T = {IN_CHANY_N32581_85,IN_CHANY_N32565_69,IN_CHANY_N32541_45}; // @[TileFull.scala 207:13]
  wire  _SBMux_C49_N23475_O_0_C_4_io_in_WIRE_1 = IN_CHANY_N32577_81; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C49_N23475_O_0_C_4_io_in_WIRE_0 = IN_CHANY_N32537_41; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C49_N23475_O_0_C_4_io_in_lo = {IN_CHANY_N32577_81,IN_CHANY_N32537_41}; // @[TileFull.scala 207:13]
  wire  _SBMux_C49_N23475_O_0_C_4_io_in_WIRE_3 = IN_CHANY_N32601_105; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C49_N23475_O_0_C_4_io_in_WIRE_2 = IN_CHANY_N32597_101; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C49_N23475_O_0_C_4_io_in_hi = {IN_CHANY_N32601_105,IN_CHANY_N32597_101}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C49_N23475_O_0_C_4_io_in_T = {IN_CHANY_N32601_105,IN_CHANY_N32597_101,IN_CHANY_N32577_81,
    IN_CHANY_N32537_41}; // @[TileFull.scala 207:13]
  wire  _SBMux_C57_N23477_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32595_99; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C57_N23477_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32563_67; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C57_N23477_O_0_C_3_io_in_hi = {IN_CHANY_N32595_99,IN_CHANY_N32563_67}; // @[TileFull.scala 207:13]
  wire  _SBMux_C57_N23477_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32499_3; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C57_N23477_O_0_C_3_io_in_T = {IN_CHANY_N32595_99,IN_CHANY_N32563_67,IN_CHANY_N32499_3}; // @[TileFull.scala 207:13]
  wire  _SBMux_C65_N23479_O_0_C_4_io_in_WIRE_1 = IN_CHANY_N32567_71; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C65_N23479_O_0_C_4_io_in_WIRE_0 = IN_CHANY_N32517_21; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C65_N23479_O_0_C_4_io_in_lo = {IN_CHANY_N32567_71,IN_CHANY_N32517_21}; // @[TileFull.scala 207:13]
  wire  _SBMux_C65_N23479_O_0_C_4_io_in_WIRE_3 = IN_CHANY_N32603_107; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C65_N23479_O_0_C_4_io_in_WIRE_2 = IN_CHANY_N32579_83; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C65_N23479_O_0_C_4_io_in_hi = {IN_CHANY_N32603_107,IN_CHANY_N32579_83}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C65_N23479_O_0_C_4_io_in_T = {IN_CHANY_N32603_107,IN_CHANY_N32579_83,IN_CHANY_N32567_71,
    IN_CHANY_N32517_21}; // @[TileFull.scala 207:13]
  wire  _SBMux_C73_N23481_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32585_89; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C73_N23481_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32565_69; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C73_N23481_O_0_C_2_io_in_T = {IN_CHANY_N32585_89,IN_CHANY_N32565_69}; // @[TileFull.scala 207:13]
  wire  _SBMux_C81_N23483_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32595_99; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C81_N23483_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32577_81; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C81_N23483_O_0_C_2_io_in_T = {IN_CHANY_N32595_99,IN_CHANY_N32577_81}; // @[TileFull.scala 207:13]
  wire  _SBMux_C3_N23497_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32593_97; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C3_N23497_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32569_73; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C3_N23497_O_0_C_3_io_in_hi = {IN_CHANY_N32593_97,IN_CHANY_N32569_73}; // @[TileFull.scala 207:13]
  wire  _SBMux_C3_N23497_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32525_29; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C3_N23497_O_0_C_3_io_in_T = {IN_CHANY_N32593_97,IN_CHANY_N32569_73,IN_CHANY_N32525_29}; // @[TileFull.scala 207:13]
  wire  _SBMux_C11_N23499_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32587_91; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C11_N23499_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32569_73; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C11_N23499_O_0_C_3_io_in_hi = {IN_CHANY_N32587_91,IN_CHANY_N32569_73}; // @[TileFull.scala 207:13]
  wire  _SBMux_C11_N23499_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32523_27; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C11_N23499_O_0_C_3_io_in_T = {IN_CHANY_N32587_91,IN_CHANY_N32569_73,IN_CHANY_N32523_27}; // @[TileFull.scala 207:13]
  wire  _SBMux_C19_N23501_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32599_103; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C19_N23501_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32571_75; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C19_N23501_O_0_C_3_io_in_hi = {IN_CHANY_N32599_103,IN_CHANY_N32571_75}; // @[TileFull.scala 207:13]
  wire  _SBMux_C19_N23501_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32515_19; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C19_N23501_O_0_C_3_io_in_T = {IN_CHANY_N32599_103,IN_CHANY_N32571_75,IN_CHANY_N32515_19}; // @[TileFull.scala 207:13]
  wire  _SBMux_C27_N23503_O_0_C_4_io_in_WIRE_1 = IN_CHANY_N32571_75; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C27_N23503_O_0_C_4_io_in_WIRE_0 = IN_CHANY_N32539_43; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C27_N23503_O_0_C_4_io_in_lo = {IN_CHANY_N32571_75,IN_CHANY_N32539_43}; // @[TileFull.scala 207:13]
  wire  _SBMux_C27_N23503_O_0_C_4_io_in_WIRE_3 = IN_CHANY_N32591_95; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C27_N23503_O_0_C_4_io_in_WIRE_2 = IN_CHANY_N32587_91; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C27_N23503_O_0_C_4_io_in_hi = {IN_CHANY_N32591_95,IN_CHANY_N32587_91}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C27_N23503_O_0_C_4_io_in_T = {IN_CHANY_N32591_95,IN_CHANY_N32587_91,IN_CHANY_N32571_75,
    IN_CHANY_N32539_43}; // @[TileFull.scala 207:13]
  wire  _SBMux_C35_N23505_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32599_103; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C35_N23505_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32575_79; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C35_N23505_O_0_C_3_io_in_hi = {IN_CHANY_N32599_103,IN_CHANY_N32575_79}; // @[TileFull.scala 207:13]
  wire  _SBMux_C35_N23505_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32507_11; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C35_N23505_O_0_C_3_io_in_T = {IN_CHANY_N32599_103,IN_CHANY_N32575_79,IN_CHANY_N32507_11}; // @[TileFull.scala 207:13]
  wire  _SBMux_C43_N23507_O_0_C_4_io_in_WIRE_1 = IN_CHANY_N32573_77; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C43_N23507_O_0_C_4_io_in_WIRE_0 = IN_CHANY_N32543_47; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C43_N23507_O_0_C_4_io_in_lo = {IN_CHANY_N32573_77,IN_CHANY_N32543_47}; // @[TileFull.scala 207:13]
  wire  _SBMux_C43_N23507_O_0_C_4_io_in_WIRE_3 = IN_CHANY_N32595_99; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C43_N23507_O_0_C_4_io_in_WIRE_2 = IN_CHANY_N32589_93; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C43_N23507_O_0_C_4_io_in_hi = {IN_CHANY_N32595_99,IN_CHANY_N32589_93}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C43_N23507_O_0_C_4_io_in_T = {IN_CHANY_N32595_99,IN_CHANY_N32589_93,IN_CHANY_N32573_77,
    IN_CHANY_N32543_47}; // @[TileFull.scala 207:13]
  wire  _SBMux_C51_N23509_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32563_67; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C51_N23509_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32553_57; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C51_N23509_O_0_C_2_io_in_T = {IN_CHANY_N32563_67,IN_CHANY_N32553_57}; // @[TileFull.scala 207:13]
  wire  _SBMux_C59_N23511_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32585_89; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C59_N23511_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32575_79; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C59_N23511_O_0_C_3_io_in_hi = {IN_CHANY_N32585_89,IN_CHANY_N32575_79}; // @[TileFull.scala 207:13]
  wire  _SBMux_C59_N23511_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32497_1; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C59_N23511_O_0_C_3_io_in_T = {IN_CHANY_N32585_89,IN_CHANY_N32575_79,IN_CHANY_N32497_1}; // @[TileFull.scala 207:13]
  wire  _SBMux_C67_N23513_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32593_97; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C67_N23513_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32575_79; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C67_N23513_O_0_C_2_io_in_T = {IN_CHANY_N32593_97,IN_CHANY_N32575_79}; // @[TileFull.scala 207:13]
  wire  _SBMux_C75_N23515_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32591_95; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C75_N23515_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32571_75; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C75_N23515_O_0_C_2_io_in_T = {IN_CHANY_N32591_95,IN_CHANY_N32571_75}; // @[TileFull.scala 207:13]
  wire  _SBMux_C83_N23517_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32603_107; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C83_N23517_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32539_43; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C83_N23517_O_0_C_2_io_in_T = {IN_CHANY_N32603_107,IN_CHANY_N32539_43}; // @[TileFull.scala 207:13]
  wire  _SBMux_C87_N23519_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32581_85; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C87_N23519_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32511_15; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C87_N23519_O_0_C_2_io_in_T = {IN_CHANY_N32581_85,IN_CHANY_N32511_15}; // @[TileFull.scala 207:13]
  wire  _SBMux_C91_N23521_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32585_89; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C91_N23521_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32497_1; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C91_N23521_O_0_C_2_io_in_T = {IN_CHANY_N32585_89,IN_CHANY_N32497_1}; // @[TileFull.scala 207:13]
  wire  _SBMux_C95_N23523_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32601_105; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C95_N23523_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32519_23; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C95_N23523_O_0_C_2_io_in_T = {IN_CHANY_N32601_105,IN_CHANY_N32519_23}; // @[TileFull.scala 207:13]
  wire  _SBMux_C99_N23525_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32579_83; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C99_N23525_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32547_51; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C99_N23525_O_0_C_2_io_in_T = {IN_CHANY_N32579_83,IN_CHANY_N32547_51}; // @[TileFull.scala 207:13]
  wire  _SBMux_C103_N23527_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32583_87; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C103_N23527_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32525_29; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C103_N23527_O_0_C_2_io_in_T = {IN_CHANY_N32583_87,IN_CHANY_N32525_29}; // @[TileFull.scala 207:13]
  wire  _SBMux_C107_N23529_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32597_101; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C107_N23529_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32517_21; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C107_N23529_O_0_C_2_io_in_T = {IN_CHANY_N32597_101,IN_CHANY_N32517_21}; // @[TileFull.scala 207:13]
  wire  _SBMux_C5_N23531_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32567_71; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C5_N23531_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32549_53; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C5_N23531_O_0_C_2_io_in_T = {IN_CHANY_N32567_71,IN_CHANY_N32549_53}; // @[TileFull.scala 207:13]
  wire  _SBMux_C13_N23533_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32577_81; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C13_N23533_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32503_7; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C13_N23533_O_0_C_2_io_in_T = {IN_CHANY_N32577_81,IN_CHANY_N32503_7}; // @[TileFull.scala 207:13]
  wire  _SBMux_C21_N23535_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32603_107; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C21_N23535_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32573_77; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C21_N23535_O_0_C_3_io_in_hi = {IN_CHANY_N32603_107,IN_CHANY_N32573_77}; // @[TileFull.scala 207:13]
  wire  _SBMux_C21_N23535_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32547_51; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C21_N23535_O_0_C_3_io_in_T = {IN_CHANY_N32603_107,IN_CHANY_N32573_77,IN_CHANY_N32547_51}; // @[TileFull.scala 207:13]
  wire  _SBMux_C29_N23537_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32579_83; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C29_N23537_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32557_61; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C29_N23537_O_0_C_2_io_in_T = {IN_CHANY_N32579_83,IN_CHANY_N32557_61}; // @[TileFull.scala 207:13]
  wire  _SBMux_C37_N23539_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32595_99; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C37_N23539_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32565_69; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C37_N23539_O_0_C_3_io_in_hi = {IN_CHANY_N32595_99,IN_CHANY_N32565_69}; // @[TileFull.scala 207:13]
  wire  _SBMux_C37_N23539_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32527_31; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C37_N23539_O_0_C_3_io_in_T = {IN_CHANY_N32595_99,IN_CHANY_N32565_69,IN_CHANY_N32527_31}; // @[TileFull.scala 207:13]
  wire  _SBMux_C45_N23541_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32569_73; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C45_N23541_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32545_49; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C45_N23541_O_0_C_2_io_in_T = {IN_CHANY_N32569_73,IN_CHANY_N32545_49}; // @[TileFull.scala 207:13]
  wire  _SBMux_C53_N23543_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32597_101; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C53_N23543_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32565_69; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C53_N23543_O_0_C_3_io_in_hi = {IN_CHANY_N32597_101,IN_CHANY_N32565_69}; // @[TileFull.scala 207:13]
  wire  _SBMux_C53_N23543_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32521_25; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C53_N23543_O_0_C_3_io_in_T = {IN_CHANY_N32597_101,IN_CHANY_N32565_69,IN_CHANY_N32521_25}; // @[TileFull.scala 207:13]
  wire  _SBMux_C61_N23545_O_0_C_3_io_in_WIRE_2 = IN_CHANY_N32581_85; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C61_N23545_O_0_C_3_io_in_WIRE_1 = IN_CHANY_N32567_71; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C61_N23545_O_0_C_3_io_in_hi = {IN_CHANY_N32581_85,IN_CHANY_N32567_71}; // @[TileFull.scala 207:13]
  wire  _SBMux_C61_N23545_O_0_C_3_io_in_WIRE_0 = IN_CHANY_N32519_23; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C61_N23545_O_0_C_3_io_in_T = {IN_CHANY_N32581_85,IN_CHANY_N32567_71,IN_CHANY_N32519_23}; // @[TileFull.scala 207:13]
  wire  _SBMux_C69_N23547_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32579_83; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C69_N23547_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32569_73; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C69_N23547_O_0_C_2_io_in_T = {IN_CHANY_N32579_83,IN_CHANY_N32569_73}; // @[TileFull.scala 207:13]
  wire  _SBMux_C77_N23549_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32587_91; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C77_N23549_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32573_77; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C77_N23549_O_0_C_2_io_in_T = {IN_CHANY_N32587_91,IN_CHANY_N32573_77}; // @[TileFull.scala 207:13]
  wire  _SBMux_C85_N23551_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32589_93; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C85_N23551_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32557_61; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C85_N23551_O_0_C_2_io_in_T = {IN_CHANY_N32589_93,IN_CHANY_N32557_61}; // @[TileFull.scala 207:13]
  wire  _SBMux_C89_N23553_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32595_99; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C89_N23553_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32537_41; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C89_N23553_O_0_C_2_io_in_T = {IN_CHANY_N32595_99,IN_CHANY_N32537_41}; // @[TileFull.scala 207:13]
  wire  _SBMux_C93_N23555_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32593_97; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C93_N23555_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32551_55; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C93_N23555_O_0_C_2_io_in_T = {IN_CHANY_N32593_97,IN_CHANY_N32551_55}; // @[TileFull.scala 207:13]
  wire  _SBMux_C97_N23557_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32587_91; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C97_N23557_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32543_47; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C97_N23557_O_0_C_2_io_in_T = {IN_CHANY_N32587_91,IN_CHANY_N32543_47}; // @[TileFull.scala 207:13]
  wire  _SBMux_C101_N23559_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32599_103; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C101_N23559_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32545_49; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C101_N23559_O_0_C_2_io_in_T = {IN_CHANY_N32599_103,IN_CHANY_N32545_49}; // @[TileFull.scala 207:13]
  wire  _SBMux_C105_N23561_O_0_C_2_io_in_WIRE_1 = IN_CHANY_N32591_95; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C105_N23561_O_0_C_2_io_in_WIRE_0 = IN_CHANY_N32561_65; // @[TileFull.scala 192:{39,39}]
  wire [1:0] _SBMux_C105_N23561_O_0_C_2_io_in_T = {IN_CHANY_N32591_95,IN_CHANY_N32561_65}; // @[TileFull.scala 207:13]
  wire  _SBMux_C0_N32496_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21952_48; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C0_N32496_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21936_32; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C0_N32496_O_2_C_3_io_in_lo = {IN_OPIN_N21952_48,IN_OPIN_N21936_32}; // @[TileFull.scala 207:13]
  wire  _SBMux_C0_N32496_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23552_88; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C0_N32496_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23496_2; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C0_N32496_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23552_88,IN_CHANX_N23496_2}; // @[TileFull.scala 207:13]
  wire  _SBMux_C0_N32496_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23482_80; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C0_N32496_O_2_C_3_io_in_hi = {IN_CHANX_N23552_88,IN_CHANX_N23496_2,IN_CHANX_N23482_80}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C0_N32496_O_2_C_3_io_in_T = {IN_CHANX_N23552_88,IN_CHANX_N23496_2,IN_CHANX_N23482_80,
    IN_OPIN_N21952_48,IN_OPIN_N21936_32}; // @[TileFull.scala 207:13]
  wire  _SBMux_C2_N32498_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21953_49; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C2_N32498_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21936_32; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C2_N32498_O_2_C_3_io_in_lo = {IN_OPIN_N21953_49,IN_OPIN_N21936_32}; // @[TileFull.scala 207:13]
  wire  _SBMux_C2_N32498_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23526_102; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C2_N32498_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23466_16; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C2_N32498_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23526_102,IN_CHANX_N23466_16}; // @[TileFull.scala 207:13]
  wire  _SBMux_C2_N32498_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23446_78; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C2_N32498_O_2_C_3_io_in_hi = {IN_CHANX_N23526_102,IN_CHANX_N23466_16,IN_CHANX_N23446_78}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C2_N32498_O_2_C_3_io_in_T = {IN_CHANX_N23526_102,IN_CHANX_N23466_16,IN_CHANX_N23446_78,
    IN_OPIN_N21953_49,IN_OPIN_N21936_32}; // @[TileFull.scala 207:13]
  wire  _SBMux_C4_N32500_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21953_49; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C4_N32500_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21937_33; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C4_N32500_O_2_C_3_io_in_lo = {IN_OPIN_N21953_49,IN_OPIN_N21937_33}; // @[TileFull.scala 207:13]
  wire  _SBMux_C4_N32500_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23548_76; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C4_N32500_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23518_86; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C4_N32500_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23548_76,IN_CHANX_N23518_86}; // @[TileFull.scala 207:13]
  wire  _SBMux_C4_N32500_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23510_58; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C4_N32500_O_2_C_3_io_in_hi = {IN_CHANX_N23548_76,IN_CHANX_N23518_86,IN_CHANX_N23510_58}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C4_N32500_O_2_C_3_io_in_T = {IN_CHANX_N23548_76,IN_CHANX_N23518_86,IN_CHANX_N23510_58,
    IN_OPIN_N21953_49,IN_OPIN_N21937_33}; // @[TileFull.scala 207:13]
  wire  _SBMux_C6_N32502_O_2_C_4_io_in_WIRE_2 = IN_CHANX_N23462_0; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C6_N32502_O_2_C_4_io_in_WIRE_1 = IN_OPIN_N21954_50; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C6_N32502_O_2_C_4_io_in_lo_hi = {IN_CHANX_N23462_0,IN_OPIN_N21954_50}; // @[TileFull.scala 207:13]
  wire  _SBMux_C6_N32502_O_2_C_4_io_in_WIRE_0 = IN_OPIN_N21937_33; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C6_N32502_O_2_C_4_io_in_lo = {IN_CHANX_N23462_0,IN_OPIN_N21954_50,IN_OPIN_N21937_33}; // @[TileFull.scala 207:13]
  wire  _SBMux_C6_N32502_O_2_C_4_io_in_WIRE_5 = IN_CHANX_N23558_100; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C6_N32502_O_2_C_4_io_in_WIRE_4 = IN_CHANX_N23554_92; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C6_N32502_O_2_C_4_io_in_hi_hi = {IN_CHANX_N23558_100,IN_CHANX_N23554_92}; // @[TileFull.scala 207:13]
  wire  _SBMux_C6_N32502_O_2_C_4_io_in_WIRE_3 = IN_CHANX_N23482_80; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C6_N32502_O_2_C_4_io_in_hi = {IN_CHANX_N23558_100,IN_CHANX_N23554_92,IN_CHANX_N23482_80}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C6_N32502_O_2_C_4_io_in_T = {IN_CHANX_N23558_100,IN_CHANX_N23554_92,IN_CHANX_N23482_80,
    IN_CHANX_N23462_0,IN_OPIN_N21954_50,IN_OPIN_N21937_33}; // @[TileFull.scala 207:13]
  wire  _SBMux_C8_N32504_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21954_50; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C8_N32504_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21938_34; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C8_N32504_O_2_C_3_io_in_lo = {IN_OPIN_N21954_50,IN_OPIN_N21938_34}; // @[TileFull.scala 207:13]
  wire  _SBMux_C8_N32504_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23532_12; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C8_N32504_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23528_106; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C8_N32504_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23532_12,IN_CHANX_N23528_106}; // @[TileFull.scala 207:13]
  wire  _SBMux_C8_N32504_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23444_70; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C8_N32504_O_2_C_3_io_in_hi = {IN_CHANX_N23532_12,IN_CHANX_N23528_106,IN_CHANX_N23444_70}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C8_N32504_O_2_C_3_io_in_T = {IN_CHANX_N23532_12,IN_CHANX_N23528_106,IN_CHANX_N23444_70,
    IN_OPIN_N21954_50,IN_OPIN_N21938_34}; // @[TileFull.scala 207:13]
  wire  _SBMux_C10_N32506_O_2_C_4_io_in_WIRE_2 = IN_CHANX_N23440_54; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C10_N32506_O_2_C_4_io_in_WIRE_1 = IN_OPIN_N21955_51; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C10_N32506_O_2_C_4_io_in_lo_hi = {IN_CHANX_N23440_54,IN_OPIN_N21955_51}; // @[TileFull.scala 207:13]
  wire  _SBMux_C10_N32506_O_2_C_4_io_in_WIRE_0 = IN_OPIN_N21938_34; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C10_N32506_O_2_C_4_io_in_lo = {IN_CHANX_N23440_54,IN_OPIN_N21955_51,IN_OPIN_N21938_34}; // @[TileFull.scala 207:13]
  wire  _SBMux_C10_N32506_O_2_C_4_io_in_WIRE_5 = IN_CHANX_N23556_96; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C10_N32506_O_2_C_4_io_in_WIRE_4 = IN_CHANX_N23550_84; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C10_N32506_O_2_C_4_io_in_hi_hi = {IN_CHANX_N23556_96,IN_CHANX_N23550_84}; // @[TileFull.scala 207:13]
  wire  _SBMux_C10_N32506_O_2_C_4_io_in_WIRE_3 = IN_CHANX_N23480_72; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C10_N32506_O_2_C_4_io_in_hi = {IN_CHANX_N23556_96,IN_CHANX_N23550_84,IN_CHANX_N23480_72}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C10_N32506_O_2_C_4_io_in_T = {IN_CHANX_N23556_96,IN_CHANX_N23550_84,IN_CHANX_N23480_72,
    IN_CHANX_N23440_54,IN_OPIN_N21955_51,IN_OPIN_N21938_34}; // @[TileFull.scala 207:13]
  wire  _SBMux_C12_N32508_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21955_51; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C12_N32508_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21939_35; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C12_N32508_O_2_C_3_io_in_lo = {IN_OPIN_N21955_51,IN_OPIN_N21939_35}; // @[TileFull.scala 207:13]
  wire  _SBMux_C12_N32508_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23546_68; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C12_N32508_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23516_82; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C12_N32508_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23546_68,IN_CHANX_N23516_82}; // @[TileFull.scala 207:13]
  wire  _SBMux_C12_N32508_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23472_40; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C12_N32508_O_2_C_3_io_in_hi = {IN_CHANX_N23546_68,IN_CHANX_N23516_82,IN_CHANX_N23472_40}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C12_N32508_O_2_C_3_io_in_T = {IN_CHANX_N23546_68,IN_CHANX_N23516_82,IN_CHANX_N23472_40,
    IN_OPIN_N21955_51,IN_OPIN_N21939_35}; // @[TileFull.scala 207:13]
  wire  _SBMux_C14_N32510_O_2_C_4_io_in_WIRE_2 = IN_CHANX_N23504_34; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C14_N32510_O_2_C_4_io_in_WIRE_1 = IN_OPIN_N21956_52; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C14_N32510_O_2_C_4_io_in_lo_hi = {IN_CHANX_N23504_34,IN_OPIN_N21956_52}; // @[TileFull.scala 207:13]
  wire  _SBMux_C14_N32510_O_2_C_4_io_in_WIRE_0 = IN_OPIN_N21939_35; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C14_N32510_O_2_C_4_io_in_lo = {IN_CHANX_N23504_34,IN_OPIN_N21956_52,IN_OPIN_N21939_35}; // @[TileFull.scala 207:13]
  wire  _SBMux_C14_N32510_O_2_C_4_io_in_WIRE_5 = IN_CHANX_N23548_76; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C14_N32510_O_2_C_4_io_in_WIRE_4 = IN_CHANX_N23522_94; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C14_N32510_O_2_C_4_io_in_hi_hi = {IN_CHANX_N23548_76,IN_CHANX_N23522_94}; // @[TileFull.scala 207:13]
  wire  _SBMux_C14_N32510_O_2_C_4_io_in_WIRE_3 = IN_CHANX_N23520_90; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C14_N32510_O_2_C_4_io_in_hi = {IN_CHANX_N23548_76,IN_CHANX_N23522_94,IN_CHANX_N23520_90}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C14_N32510_O_2_C_4_io_in_T = {IN_CHANX_N23548_76,IN_CHANX_N23522_94,IN_CHANX_N23520_90,
    IN_CHANX_N23504_34,IN_OPIN_N21956_52,IN_OPIN_N21939_35}; // @[TileFull.scala 207:13]
  wire  _SBMux_C16_N32512_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21956_52; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C16_N32512_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21940_36; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C16_N32512_O_2_C_3_io_in_lo = {IN_OPIN_N21956_52,IN_OPIN_N21940_36}; // @[TileFull.scala 207:13]
  wire  _SBMux_C16_N32512_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23548_76; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C16_N32512_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23528_106; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C16_N32512_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23548_76,IN_CHANX_N23528_106}; // @[TileFull.scala 207:13]
  wire  _SBMux_C16_N32512_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23438_46; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C16_N32512_O_2_C_3_io_in_hi = {IN_CHANX_N23548_76,IN_CHANX_N23528_106,IN_CHANX_N23438_46}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C16_N32512_O_2_C_3_io_in_T = {IN_CHANX_N23548_76,IN_CHANX_N23528_106,IN_CHANX_N23438_46,
    IN_OPIN_N21956_52,IN_OPIN_N21940_36}; // @[TileFull.scala 207:13]
  wire  _SBMux_C18_N32514_O_2_C_4_io_in_WIRE_2 = IN_CHANX_N23480_72; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C18_N32514_O_2_C_4_io_in_WIRE_1 = IN_OPIN_N21957_53; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C18_N32514_O_2_C_4_io_in_lo_hi = {IN_CHANX_N23480_72,IN_OPIN_N21957_53}; // @[TileFull.scala 207:13]
  wire  _SBMux_C18_N32514_O_2_C_4_io_in_WIRE_0 = IN_OPIN_N21940_36; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C18_N32514_O_2_C_4_io_in_lo = {IN_CHANX_N23480_72,IN_OPIN_N21957_53,IN_OPIN_N21940_36}; // @[TileFull.scala 207:13]
  wire  _SBMux_C18_N32514_O_2_C_4_io_in_WIRE_5 = IN_CHANX_N23552_88; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C18_N32514_O_2_C_4_io_in_WIRE_4 = IN_CHANX_N23540_44; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C18_N32514_O_2_C_4_io_in_hi_hi = {IN_CHANX_N23552_88,IN_CHANX_N23540_44}; // @[TileFull.scala 207:13]
  wire  _SBMux_C18_N32514_O_2_C_4_io_in_WIRE_3 = IN_CHANX_N23528_106; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C18_N32514_O_2_C_4_io_in_hi = {IN_CHANX_N23552_88,IN_CHANX_N23540_44,IN_CHANX_N23528_106}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C18_N32514_O_2_C_4_io_in_T = {IN_CHANX_N23552_88,IN_CHANX_N23540_44,IN_CHANX_N23528_106,
    IN_CHANX_N23480_72,IN_OPIN_N21957_53,IN_OPIN_N21940_36}; // @[TileFull.scala 207:13]
  wire  _SBMux_C20_N32516_O_2_C_4_io_in_WIRE_2 = IN_CHANX_N23482_80; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C20_N32516_O_2_C_4_io_in_WIRE_1 = IN_OPIN_N21957_53; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C20_N32516_O_2_C_4_io_in_lo_hi = {IN_CHANX_N23482_80,IN_OPIN_N21957_53}; // @[TileFull.scala 207:13]
  wire  _SBMux_C20_N32516_O_2_C_4_io_in_WIRE_0 = IN_OPIN_N21941_37; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C20_N32516_O_2_C_4_io_in_lo = {IN_CHANX_N23482_80,IN_OPIN_N21957_53,IN_OPIN_N21941_37}; // @[TileFull.scala 207:13]
  wire  _SBMux_C20_N32516_O_2_C_4_io_in_WIRE_5 = IN_CHANX_N23560_104; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C20_N32516_O_2_C_4_io_in_WIRE_4 = IN_CHANX_N23534_20; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C20_N32516_O_2_C_4_io_in_hi_hi = {IN_CHANX_N23560_104,IN_CHANX_N23534_20}; // @[TileFull.scala 207:13]
  wire  _SBMux_C20_N32516_O_2_C_4_io_in_WIRE_3 = IN_CHANX_N23516_82; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C20_N32516_O_2_C_4_io_in_hi = {IN_CHANX_N23560_104,IN_CHANX_N23534_20,IN_CHANX_N23516_82}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C20_N32516_O_2_C_4_io_in_T = {IN_CHANX_N23560_104,IN_CHANX_N23534_20,IN_CHANX_N23516_82,
    IN_CHANX_N23482_80,IN_OPIN_N21957_53,IN_OPIN_N21941_37}; // @[TileFull.scala 207:13]
  wire  _SBMux_C22_N32518_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21958_54; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C22_N32518_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21941_37; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C22_N32518_O_2_C_3_io_in_lo = {IN_OPIN_N21958_54,IN_OPIN_N21941_37}; // @[TileFull.scala 207:13]
  wire  _SBMux_C22_N32518_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23546_68; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C22_N32518_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23520_90; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C22_N32518_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23546_68,IN_CHANX_N23520_90}; // @[TileFull.scala 207:13]
  wire  _SBMux_C22_N32518_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23476_56; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C22_N32518_O_2_C_3_io_in_hi = {IN_CHANX_N23546_68,IN_CHANX_N23520_90,IN_CHANX_N23476_56}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C22_N32518_O_2_C_3_io_in_T = {IN_CHANX_N23546_68,IN_CHANX_N23520_90,IN_CHANX_N23476_56,
    IN_OPIN_N21958_54,IN_OPIN_N21941_37}; // @[TileFull.scala 207:13]
  wire  _SBMux_C24_N32520_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21958_54; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C24_N32520_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21942_38; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C24_N32520_O_2_C_2_io_in_lo = {IN_OPIN_N21958_54,IN_OPIN_N21942_38}; // @[TileFull.scala 207:13]
  wire  _SBMux_C24_N32520_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23548_76; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C24_N32520_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23432_22; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C24_N32520_O_2_C_2_io_in_hi = {IN_CHANX_N23548_76,IN_CHANX_N23432_22}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C24_N32520_O_2_C_2_io_in_T = {IN_CHANX_N23548_76,IN_CHANX_N23432_22,IN_OPIN_N21958_54,
    IN_OPIN_N21942_38}; // @[TileFull.scala 207:13]
  wire  _SBMux_C26_N32522_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21959_55; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C26_N32522_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21942_38; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C26_N32522_O_2_C_3_io_in_lo = {IN_OPIN_N21959_55,IN_OPIN_N21942_38}; // @[TileFull.scala 207:13]
  wire  _SBMux_C26_N32522_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23550_84; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C26_N32522_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23470_32; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C26_N32522_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23550_84,IN_CHANX_N23470_32}; // @[TileFull.scala 207:13]
  wire  _SBMux_C26_N32522_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23446_78; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C26_N32522_O_2_C_3_io_in_hi = {IN_CHANX_N23550_84,IN_CHANX_N23470_32,IN_CHANX_N23446_78}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C26_N32522_O_2_C_3_io_in_T = {IN_CHANX_N23550_84,IN_CHANX_N23470_32,IN_CHANX_N23446_78,
    IN_OPIN_N21959_55,IN_OPIN_N21942_38}; // @[TileFull.scala 207:13]
  wire  _SBMux_C28_N32524_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21959_55; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C28_N32524_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21943_39; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C28_N32524_O_2_C_2_io_in_lo = {IN_OPIN_N21959_55,IN_OPIN_N21943_39}; // @[TileFull.scala 207:13]
  wire  _SBMux_C28_N32524_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23514_74; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C28_N32524_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23498_10; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C28_N32524_O_2_C_2_io_in_hi = {IN_CHANX_N23514_74,IN_CHANX_N23498_10}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C28_N32524_O_2_C_2_io_in_T = {IN_CHANX_N23514_74,IN_CHANX_N23498_10,IN_OPIN_N21959_55,
    IN_OPIN_N21943_39}; // @[TileFull.scala 207:13]
  wire  _SBMux_C30_N32526_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21960_56; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C30_N32526_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21943_39; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C30_N32526_O_2_C_2_io_in_lo = {IN_OPIN_N21960_56,IN_OPIN_N21943_39}; // @[TileFull.scala 207:13]
  wire  _SBMux_C30_N32526_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23536_28; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C30_N32526_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23444_70; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C30_N32526_O_2_C_2_io_in_hi = {IN_CHANX_N23536_28,IN_CHANX_N23444_70}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C30_N32526_O_2_C_2_io_in_T = {IN_CHANX_N23536_28,IN_CHANX_N23444_70,IN_OPIN_N21960_56,
    IN_OPIN_N21943_39}; // @[TileFull.scala 207:13]
  wire  _SBMux_C32_N32528_O_2_C_4_io_in_WIRE_2 = IN_CHANX_N23508_50; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C32_N32528_O_2_C_4_io_in_WIRE_1 = IN_OPIN_N21960_56; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C32_N32528_O_2_C_4_io_in_lo_hi = {IN_CHANX_N23508_50,IN_OPIN_N21960_56}; // @[TileFull.scala 207:13]
  wire  _SBMux_C32_N32528_O_2_C_4_io_in_WIRE_0 = IN_OPIN_N21944_40; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C32_N32528_O_2_C_4_io_in_lo = {IN_CHANX_N23508_50,IN_OPIN_N21960_56,IN_OPIN_N21944_40}; // @[TileFull.scala 207:13]
  wire  _SBMux_C32_N32528_O_2_C_4_io_in_WIRE_5 = IN_CHANX_N23524_98; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C32_N32528_O_2_C_4_io_in_WIRE_4 = IN_CHANX_N23518_86; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C32_N32528_O_2_C_4_io_in_hi_hi = {IN_CHANX_N23524_98,IN_CHANX_N23518_86}; // @[TileFull.scala 207:13]
  wire  _SBMux_C32_N32528_O_2_C_4_io_in_WIRE_3 = IN_CHANX_N23512_66; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C32_N32528_O_2_C_4_io_in_hi = {IN_CHANX_N23524_98,IN_CHANX_N23518_86,IN_CHANX_N23512_66}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C32_N32528_O_2_C_4_io_in_T = {IN_CHANX_N23524_98,IN_CHANX_N23518_86,IN_CHANX_N23512_66,
    IN_CHANX_N23508_50,IN_OPIN_N21960_56,IN_OPIN_N21944_40}; // @[TileFull.scala 207:13]
  wire  _SBMux_C34_N32530_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21961_57; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C34_N32530_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21944_40; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C34_N32530_O_2_C_3_io_in_lo = {IN_OPIN_N21961_57,IN_OPIN_N21944_40}; // @[TileFull.scala 207:13]
  wire  _SBMux_C34_N32530_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23554_92; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C34_N32530_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23542_52; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C34_N32530_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23554_92,IN_CHANX_N23542_52}; // @[TileFull.scala 207:13]
  wire  _SBMux_C34_N32530_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23480_72; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C34_N32530_O_2_C_3_io_in_hi = {IN_CHANX_N23554_92,IN_CHANX_N23542_52,IN_CHANX_N23480_72}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C34_N32530_O_2_C_3_io_in_T = {IN_CHANX_N23554_92,IN_CHANX_N23542_52,IN_CHANX_N23480_72,
    IN_OPIN_N21961_57,IN_OPIN_N21944_40}; // @[TileFull.scala 207:13]
  wire  _SBMux_C36_N32532_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21961_57; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C36_N32532_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21945_41; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C36_N32532_O_2_C_3_io_in_lo = {IN_OPIN_N21961_57,IN_OPIN_N21945_41}; // @[TileFull.scala 207:13]
  wire  _SBMux_C36_N32532_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23538_36; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C36_N32532_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23526_102; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C36_N32532_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23538_36,IN_CHANX_N23526_102}; // @[TileFull.scala 207:13]
  wire  _SBMux_C36_N32532_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23480_72; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C36_N32532_O_2_C_3_io_in_hi = {IN_CHANX_N23538_36,IN_CHANX_N23526_102,IN_CHANX_N23480_72}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C36_N32532_O_2_C_3_io_in_T = {IN_CHANX_N23538_36,IN_CHANX_N23526_102,IN_CHANX_N23480_72,
    IN_OPIN_N21961_57,IN_OPIN_N21945_41}; // @[TileFull.scala 207:13]
  wire  _SBMux_C38_N32534_O_2_C_4_io_in_WIRE_2 = IN_CHANX_N23434_30; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C38_N32534_O_2_C_4_io_in_WIRE_1 = IN_OPIN_N21962_58; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C38_N32534_O_2_C_4_io_in_lo_hi = {IN_CHANX_N23434_30,IN_OPIN_N21962_58}; // @[TileFull.scala 207:13]
  wire  _SBMux_C38_N32534_O_2_C_4_io_in_WIRE_0 = IN_OPIN_N21945_41; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C38_N32534_O_2_C_4_io_in_lo = {IN_CHANX_N23434_30,IN_OPIN_N21962_58,IN_OPIN_N21945_41}; // @[TileFull.scala 207:13]
  wire  _SBMux_C38_N32534_O_2_C_4_io_in_WIRE_5 = IN_CHANX_N23560_104; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C38_N32534_O_2_C_4_io_in_WIRE_4 = IN_CHANX_N23514_74; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C38_N32534_O_2_C_4_io_in_hi_hi = {IN_CHANX_N23560_104,IN_CHANX_N23514_74}; // @[TileFull.scala 207:13]
  wire  _SBMux_C38_N32534_O_2_C_4_io_in_WIRE_3 = IN_CHANX_N23512_66; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C38_N32534_O_2_C_4_io_in_hi = {IN_CHANX_N23560_104,IN_CHANX_N23514_74,IN_CHANX_N23512_66}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C38_N32534_O_2_C_4_io_in_T = {IN_CHANX_N23560_104,IN_CHANX_N23514_74,IN_CHANX_N23512_66,
    IN_CHANX_N23434_30,IN_OPIN_N21962_58,IN_OPIN_N21945_41}; // @[TileFull.scala 207:13]
  wire  _SBMux_C40_N32536_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21962_58; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C40_N32536_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21946_42; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C40_N32536_O_2_C_2_io_in_lo = {IN_OPIN_N21962_58,IN_OPIN_N21946_42}; // @[TileFull.scala 207:13]
  wire  _SBMux_C40_N32536_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23526_102; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C40_N32536_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23506_42; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C40_N32536_O_2_C_2_io_in_hi = {IN_CHANX_N23526_102,IN_CHANX_N23506_42}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C40_N32536_O_2_C_2_io_in_T = {IN_CHANX_N23526_102,IN_CHANX_N23506_42,IN_OPIN_N21962_58,
    IN_OPIN_N21946_42}; // @[TileFull.scala 207:13]
  wire  _SBMux_C42_N32538_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21963_59; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C42_N32538_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21946_42; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C42_N32538_O_2_C_3_io_in_lo = {IN_OPIN_N21963_59,IN_OPIN_N21946_42}; // @[TileFull.scala 207:13]
  wire  _SBMux_C42_N32538_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23558_100; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C42_N32538_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23446_78; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C42_N32538_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23558_100,IN_CHANX_N23446_78}; // @[TileFull.scala 207:13]
  wire  _SBMux_C42_N32538_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23442_62; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C42_N32538_O_2_C_3_io_in_hi = {IN_CHANX_N23558_100,IN_CHANX_N23446_78,IN_CHANX_N23442_62}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C42_N32538_O_2_C_3_io_in_T = {IN_CHANX_N23558_100,IN_CHANX_N23446_78,IN_CHANX_N23442_62,
    IN_OPIN_N21963_59,IN_OPIN_N21946_42}; // @[TileFull.scala 207:13]
  wire  _SBMux_C44_N32540_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21963_59; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C44_N32540_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21947_43; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C44_N32540_O_2_C_3_io_in_lo = {IN_OPIN_N21963_59,IN_OPIN_N21947_43}; // @[TileFull.scala 207:13]
  wire  _SBMux_C44_N32540_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23520_90; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C44_N32540_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23512_66; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C44_N32540_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23520_90,IN_CHANX_N23512_66}; // @[TileFull.scala 207:13]
  wire  _SBMux_C44_N32540_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23436_38; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C44_N32540_O_2_C_3_io_in_hi = {IN_CHANX_N23520_90,IN_CHANX_N23512_66,IN_CHANX_N23436_38}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C44_N32540_O_2_C_3_io_in_T = {IN_CHANX_N23520_90,IN_CHANX_N23512_66,IN_CHANX_N23436_38,
    IN_OPIN_N21963_59,IN_OPIN_N21947_43}; // @[TileFull.scala 207:13]
  wire  _SBMux_C46_N32542_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21964_60; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C46_N32542_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21947_43; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C46_N32542_O_2_C_3_io_in_lo = {IN_OPIN_N21964_60,IN_OPIN_N21947_43}; // @[TileFull.scala 207:13]
  wire  _SBMux_C46_N32542_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23556_96; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C46_N32542_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23546_68; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C46_N32542_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23556_96,IN_CHANX_N23546_68}; // @[TileFull.scala 207:13]
  wire  _SBMux_C46_N32542_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23530_4; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C46_N32542_O_2_C_3_io_in_hi = {IN_CHANX_N23556_96,IN_CHANX_N23546_68,IN_CHANX_N23530_4}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C46_N32542_O_2_C_3_io_in_T = {IN_CHANX_N23556_96,IN_CHANX_N23546_68,IN_CHANX_N23530_4,
    IN_OPIN_N21964_60,IN_OPIN_N21947_43}; // @[TileFull.scala 207:13]
  wire  _SBMux_C48_N32544_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21964_60; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C48_N32544_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21948_44; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C48_N32544_O_2_C_3_io_in_lo = {IN_OPIN_N21964_60,IN_OPIN_N21948_44}; // @[TileFull.scala 207:13]
  wire  _SBMux_C48_N32544_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23554_92; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C48_N32544_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23512_66; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C48_N32544_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23554_92,IN_CHANX_N23512_66}; // @[TileFull.scala 207:13]
  wire  _SBMux_C48_N32544_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23464_8; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C48_N32544_O_2_C_3_io_in_hi = {IN_CHANX_N23554_92,IN_CHANX_N23512_66,IN_CHANX_N23464_8}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C48_N32544_O_2_C_3_io_in_T = {IN_CHANX_N23554_92,IN_CHANX_N23512_66,IN_CHANX_N23464_8,
    IN_OPIN_N21964_60,IN_OPIN_N21948_44}; // @[TileFull.scala 207:13]
  wire  _SBMux_C50_N32546_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21965_61; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C50_N32546_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21948_44; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C50_N32546_O_2_C_3_io_in_lo = {IN_OPIN_N21965_61,IN_OPIN_N21948_44}; // @[TileFull.scala 207:13]
  wire  _SBMux_C50_N32546_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23518_86; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C50_N32546_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23478_64; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C50_N32546_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23518_86,IN_CHANX_N23478_64}; // @[TileFull.scala 207:13]
  wire  _SBMux_C50_N32546_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23446_78; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C50_N32546_O_2_C_3_io_in_hi = {IN_CHANX_N23518_86,IN_CHANX_N23478_64,IN_CHANX_N23446_78}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C50_N32546_O_2_C_3_io_in_T = {IN_CHANX_N23518_86,IN_CHANX_N23478_64,IN_CHANX_N23446_78,
    IN_OPIN_N21965_61,IN_OPIN_N21948_44}; // @[TileFull.scala 207:13]
  wire  _SBMux_C52_N32548_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21965_61; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C52_N32548_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21949_45; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C52_N32548_O_2_C_3_io_in_lo = {IN_OPIN_N21965_61,IN_OPIN_N21949_45}; // @[TileFull.scala 207:13]
  wire  _SBMux_C52_N32548_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23522_94; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C52_N32548_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23500_18; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C52_N32548_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23522_94,IN_CHANX_N23500_18}; // @[TileFull.scala 207:13]
  wire  _SBMux_C52_N32548_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23444_70; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C52_N32548_O_2_C_3_io_in_hi = {IN_CHANX_N23522_94,IN_CHANX_N23500_18,IN_CHANX_N23444_70}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C52_N32548_O_2_C_3_io_in_T = {IN_CHANX_N23522_94,IN_CHANX_N23500_18,IN_CHANX_N23444_70,
    IN_OPIN_N21965_61,IN_OPIN_N21949_45}; // @[TileFull.scala 207:13]
  wire  _SBMux_C54_N32550_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21966_62; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C54_N32550_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21949_45; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C54_N32550_O_2_C_2_io_in_lo = {IN_OPIN_N21966_62,IN_OPIN_N21949_45}; // @[TileFull.scala 207:13]
  wire  _SBMux_C54_N32550_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23546_68; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C54_N32550_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23430_14; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C54_N32550_O_2_C_2_io_in_hi = {IN_CHANX_N23546_68,IN_CHANX_N23430_14}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C54_N32550_O_2_C_2_io_in_T = {IN_CHANX_N23546_68,IN_CHANX_N23430_14,IN_OPIN_N21966_62,
    IN_OPIN_N21949_45}; // @[TileFull.scala 207:13]
  wire  _SBMux_C56_N32552_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21966_62; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C56_N32552_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21950_46; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C56_N32552_O_2_C_3_io_in_lo = {IN_OPIN_N21966_62,IN_OPIN_N21950_46}; // @[TileFull.scala 207:13]
  wire  _SBMux_C56_N32552_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23550_84; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C56_N32552_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23482_80; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C56_N32552_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23550_84,IN_CHANX_N23482_80}; // @[TileFull.scala 207:13]
  wire  _SBMux_C56_N32552_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23474_48; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C56_N32552_O_2_C_3_io_in_hi = {IN_CHANX_N23550_84,IN_CHANX_N23482_80,IN_CHANX_N23474_48}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C56_N32552_O_2_C_3_io_in_T = {IN_CHANX_N23550_84,IN_CHANX_N23482_80,IN_CHANX_N23474_48,
    IN_OPIN_N21966_62,IN_OPIN_N21950_46}; // @[TileFull.scala 207:13]
  wire  _SBMux_C58_N32554_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21967_63; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C58_N32554_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21950_46; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C58_N32554_O_2_C_2_io_in_lo = {IN_OPIN_N21967_63,IN_OPIN_N21950_46}; // @[TileFull.scala 207:13]
  wire  _SBMux_C58_N32554_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23468_24; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C58_N32554_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23444_70; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C58_N32554_O_2_C_2_io_in_hi = {IN_CHANX_N23468_24,IN_CHANX_N23444_70}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C58_N32554_O_2_C_2_io_in_T = {IN_CHANX_N23468_24,IN_CHANX_N23444_70,IN_OPIN_N21967_63,
    IN_OPIN_N21950_46}; // @[TileFull.scala 207:13]
  wire  _SBMux_C60_N32556_O_2_C_3_io_in_WIRE_1 = IN_OPIN_N21967_63; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C60_N32556_O_2_C_3_io_in_WIRE_0 = IN_OPIN_N21951_47; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C60_N32556_O_2_C_3_io_in_lo = {IN_OPIN_N21967_63,IN_OPIN_N21951_47}; // @[TileFull.scala 207:13]
  wire  _SBMux_C60_N32556_O_2_C_3_io_in_WIRE_4 = IN_CHANX_N23544_60; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C60_N32556_O_2_C_3_io_in_WIRE_3 = IN_CHANX_N23524_98; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C60_N32556_O_2_C_3_io_in_hi_hi = {IN_CHANX_N23544_60,IN_CHANX_N23524_98}; // @[TileFull.scala 207:13]
  wire  _SBMux_C60_N32556_O_2_C_3_io_in_WIRE_2 = IN_CHANX_N23514_74; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C60_N32556_O_2_C_3_io_in_hi = {IN_CHANX_N23544_60,IN_CHANX_N23524_98,IN_CHANX_N23514_74}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C60_N32556_O_2_C_3_io_in_T = {IN_CHANX_N23544_60,IN_CHANX_N23524_98,IN_CHANX_N23514_74,
    IN_OPIN_N21967_63,IN_OPIN_N21951_47}; // @[TileFull.scala 207:13]
  wire  _SBMux_C62_N32558_O_1_C_3_io_in_WIRE_1 = IN_CHANX_N23428_6; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C62_N32558_O_1_C_3_io_in_WIRE_0 = IN_OPIN_N21951_47; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C62_N32558_O_1_C_3_io_in_lo = {IN_CHANX_N23428_6,IN_OPIN_N21951_47}; // @[TileFull.scala 207:13]
  wire  _SBMux_C62_N32558_O_1_C_3_io_in_WIRE_3 = IN_CHANX_N23516_82; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C62_N32558_O_1_C_3_io_in_WIRE_2 = IN_CHANX_N23512_66; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C62_N32558_O_1_C_3_io_in_hi = {IN_CHANX_N23516_82,IN_CHANX_N23512_66}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C62_N32558_O_1_C_3_io_in_T = {IN_CHANX_N23516_82,IN_CHANX_N23512_66,IN_CHANX_N23428_6,
    IN_OPIN_N21951_47}; // @[TileFull.scala 207:13]
  wire  _SBMux_C64_N32560_O_1_C_2_io_in_WIRE_2 = IN_CHANX_N23514_74; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C64_N32560_O_1_C_2_io_in_WIRE_1 = IN_CHANX_N23502_26; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C64_N32560_O_1_C_2_io_in_hi = {IN_CHANX_N23514_74,IN_CHANX_N23502_26}; // @[TileFull.scala 207:13]
  wire  _SBMux_C64_N32560_O_1_C_2_io_in_WIRE_0 = IN_OPIN_N21952_48; // @[TileFull.scala 192:{39,39}]
  wire [2:0] _SBMux_C64_N32560_O_1_C_2_io_in_T = {IN_CHANX_N23514_74,IN_CHANX_N23502_26,IN_OPIN_N21952_48}; // @[TileFull.scala 207:13]
  wire  _SBMux_C66_N32562_O_4_C_2_io_in_WIRE_2 = IN_OPIN_N21952_48; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C66_N32562_O_4_C_2_io_in_WIRE_1 = IN_OPIN_N21944_40; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C66_N32562_O_4_C_2_io_in_lo_hi = {IN_OPIN_N21952_48,IN_OPIN_N21944_40}; // @[TileFull.scala 207:13]
  wire  _SBMux_C66_N32562_O_4_C_2_io_in_WIRE_0 = IN_OPIN_N21936_32; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C66_N32562_O_4_C_2_io_in_lo = {IN_OPIN_N21952_48,IN_OPIN_N21944_40,IN_OPIN_N21936_32}; // @[TileFull.scala 207:13]
  wire  _SBMux_C66_N32562_O_4_C_2_io_in_WIRE_5 = IN_CHANX_N23552_88; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C66_N32562_O_4_C_2_io_in_WIRE_4 = IN_CHANX_N23512_66; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C66_N32562_O_4_C_2_io_in_hi_hi = {IN_CHANX_N23552_88,IN_CHANX_N23512_66}; // @[TileFull.scala 207:13]
  wire  _SBMux_C66_N32562_O_4_C_2_io_in_WIRE_3 = IN_OPIN_N21960_56; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C66_N32562_O_4_C_2_io_in_hi = {IN_CHANX_N23552_88,IN_CHANX_N23512_66,IN_OPIN_N21960_56}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C66_N32562_O_4_C_2_io_in_T = {IN_CHANX_N23552_88,IN_CHANX_N23512_66,IN_OPIN_N21960_56,
    IN_OPIN_N21952_48,IN_OPIN_N21944_40,IN_OPIN_N21936_32}; // @[TileFull.scala 207:13]
  wire  _SBMux_C68_N32564_O_4_C_2_io_in_WIRE_2 = IN_OPIN_N21953_49; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C68_N32564_O_4_C_2_io_in_WIRE_1 = IN_OPIN_N21945_41; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C68_N32564_O_4_C_2_io_in_lo_hi = {IN_OPIN_N21953_49,IN_OPIN_N21945_41}; // @[TileFull.scala 207:13]
  wire  _SBMux_C68_N32564_O_4_C_2_io_in_WIRE_0 = IN_OPIN_N21937_33; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C68_N32564_O_4_C_2_io_in_lo = {IN_OPIN_N21953_49,IN_OPIN_N21945_41,IN_OPIN_N21937_33}; // @[TileFull.scala 207:13]
  wire  _SBMux_C68_N32564_O_4_C_2_io_in_WIRE_5 = IN_CHANX_N23560_104; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C68_N32564_O_4_C_2_io_in_WIRE_4 = IN_CHANX_N23548_76; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C68_N32564_O_4_C_2_io_in_hi_hi = {IN_CHANX_N23560_104,IN_CHANX_N23548_76}; // @[TileFull.scala 207:13]
  wire  _SBMux_C68_N32564_O_4_C_2_io_in_WIRE_3 = IN_OPIN_N21961_57; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C68_N32564_O_4_C_2_io_in_hi = {IN_CHANX_N23560_104,IN_CHANX_N23548_76,IN_OPIN_N21961_57}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C68_N32564_O_4_C_2_io_in_T = {IN_CHANX_N23560_104,IN_CHANX_N23548_76,IN_OPIN_N21961_57,
    IN_OPIN_N21953_49,IN_OPIN_N21945_41,IN_OPIN_N21937_33}; // @[TileFull.scala 207:13]
  wire  _SBMux_C70_N32566_O_4_C_2_io_in_WIRE_2 = IN_OPIN_N21954_50; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C70_N32566_O_4_C_2_io_in_WIRE_1 = IN_OPIN_N21946_42; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C70_N32566_O_4_C_2_io_in_lo_hi = {IN_OPIN_N21954_50,IN_OPIN_N21946_42}; // @[TileFull.scala 207:13]
  wire  _SBMux_C70_N32566_O_4_C_2_io_in_WIRE_0 = IN_OPIN_N21938_34; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C70_N32566_O_4_C_2_io_in_lo = {IN_OPIN_N21954_50,IN_OPIN_N21946_42,IN_OPIN_N21938_34}; // @[TileFull.scala 207:13]
  wire  _SBMux_C70_N32566_O_4_C_2_io_in_WIRE_5 = IN_CHANX_N23526_102; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C70_N32566_O_4_C_2_io_in_WIRE_4 = IN_CHANX_N23480_72; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C70_N32566_O_4_C_2_io_in_hi_hi = {IN_CHANX_N23526_102,IN_CHANX_N23480_72}; // @[TileFull.scala 207:13]
  wire  _SBMux_C70_N32566_O_4_C_2_io_in_WIRE_3 = IN_OPIN_N21962_58; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C70_N32566_O_4_C_2_io_in_hi = {IN_CHANX_N23526_102,IN_CHANX_N23480_72,IN_OPIN_N21962_58}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C70_N32566_O_4_C_2_io_in_T = {IN_CHANX_N23526_102,IN_CHANX_N23480_72,IN_OPIN_N21962_58,
    IN_OPIN_N21954_50,IN_OPIN_N21946_42,IN_OPIN_N21938_34}; // @[TileFull.scala 207:13]
  wire  _SBMux_C72_N32568_O_4_C_2_io_in_WIRE_2 = IN_OPIN_N21955_51; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C72_N32568_O_4_C_2_io_in_WIRE_1 = IN_OPIN_N21947_43; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C72_N32568_O_4_C_2_io_in_lo_hi = {IN_OPIN_N21955_51,IN_OPIN_N21947_43}; // @[TileFull.scala 207:13]
  wire  _SBMux_C72_N32568_O_4_C_2_io_in_WIRE_0 = IN_OPIN_N21939_35; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C72_N32568_O_4_C_2_io_in_lo = {IN_OPIN_N21955_51,IN_OPIN_N21947_43,IN_OPIN_N21939_35}; // @[TileFull.scala 207:13]
  wire  _SBMux_C72_N32568_O_4_C_2_io_in_WIRE_5 = IN_CHANX_N23558_100; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C72_N32568_O_4_C_2_io_in_WIRE_4 = IN_CHANX_N23546_68; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C72_N32568_O_4_C_2_io_in_hi_hi = {IN_CHANX_N23558_100,IN_CHANX_N23546_68}; // @[TileFull.scala 207:13]
  wire  _SBMux_C72_N32568_O_4_C_2_io_in_WIRE_3 = IN_OPIN_N21963_59; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C72_N32568_O_4_C_2_io_in_hi = {IN_CHANX_N23558_100,IN_CHANX_N23546_68,IN_OPIN_N21963_59}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C72_N32568_O_4_C_2_io_in_T = {IN_CHANX_N23558_100,IN_CHANX_N23546_68,IN_OPIN_N21963_59,
    IN_OPIN_N21955_51,IN_OPIN_N21947_43,IN_OPIN_N21939_35}; // @[TileFull.scala 207:13]
  wire  _SBMux_C74_N32570_O_4_C_2_io_in_WIRE_2 = IN_OPIN_N21956_52; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C74_N32570_O_4_C_2_io_in_WIRE_1 = IN_OPIN_N21948_44; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C74_N32570_O_4_C_2_io_in_lo_hi = {IN_OPIN_N21956_52,IN_OPIN_N21948_44}; // @[TileFull.scala 207:13]
  wire  _SBMux_C74_N32570_O_4_C_2_io_in_WIRE_0 = IN_OPIN_N21940_36; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C74_N32570_O_4_C_2_io_in_lo = {IN_OPIN_N21956_52,IN_OPIN_N21948_44,IN_OPIN_N21940_36}; // @[TileFull.scala 207:13]
  wire  _SBMux_C74_N32570_O_4_C_2_io_in_WIRE_5 = IN_CHANX_N23524_98; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C74_N32570_O_4_C_2_io_in_WIRE_4 = IN_CHANX_N23482_80; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C74_N32570_O_4_C_2_io_in_hi_hi = {IN_CHANX_N23524_98,IN_CHANX_N23482_80}; // @[TileFull.scala 207:13]
  wire  _SBMux_C74_N32570_O_4_C_2_io_in_WIRE_3 = IN_OPIN_N21964_60; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C74_N32570_O_4_C_2_io_in_hi = {IN_CHANX_N23524_98,IN_CHANX_N23482_80,IN_OPIN_N21964_60}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C74_N32570_O_4_C_2_io_in_T = {IN_CHANX_N23524_98,IN_CHANX_N23482_80,IN_OPIN_N21964_60,
    IN_OPIN_N21956_52,IN_OPIN_N21948_44,IN_OPIN_N21940_36}; // @[TileFull.scala 207:13]
  wire  _SBMux_C76_N32572_O_4_C_2_io_in_WIRE_2 = IN_OPIN_N21957_53; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C76_N32572_O_4_C_2_io_in_WIRE_1 = IN_OPIN_N21949_45; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C76_N32572_O_4_C_2_io_in_lo_hi = {IN_OPIN_N21957_53,IN_OPIN_N21949_45}; // @[TileFull.scala 207:13]
  wire  _SBMux_C76_N32572_O_4_C_2_io_in_WIRE_0 = IN_OPIN_N21941_37; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C76_N32572_O_4_C_2_io_in_lo = {IN_OPIN_N21957_53,IN_OPIN_N21949_45,IN_OPIN_N21941_37}; // @[TileFull.scala 207:13]
  wire  _SBMux_C76_N32572_O_4_C_2_io_in_WIRE_5 = IN_CHANX_N23550_84; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C76_N32572_O_4_C_2_io_in_WIRE_4 = IN_CHANX_N23444_70; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C76_N32572_O_4_C_2_io_in_hi_hi = {IN_CHANX_N23550_84,IN_CHANX_N23444_70}; // @[TileFull.scala 207:13]
  wire  _SBMux_C76_N32572_O_4_C_2_io_in_WIRE_3 = IN_OPIN_N21965_61; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C76_N32572_O_4_C_2_io_in_hi = {IN_CHANX_N23550_84,IN_CHANX_N23444_70,IN_OPIN_N21965_61}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C76_N32572_O_4_C_2_io_in_T = {IN_CHANX_N23550_84,IN_CHANX_N23444_70,IN_OPIN_N21965_61,
    IN_OPIN_N21957_53,IN_OPIN_N21949_45,IN_OPIN_N21941_37}; // @[TileFull.scala 207:13]
  wire  _SBMux_C78_N32574_O_4_C_2_io_in_WIRE_2 = IN_OPIN_N21958_54; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C78_N32574_O_4_C_2_io_in_WIRE_1 = IN_OPIN_N21950_46; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C78_N32574_O_4_C_2_io_in_lo_hi = {IN_OPIN_N21958_54,IN_OPIN_N21950_46}; // @[TileFull.scala 207:13]
  wire  _SBMux_C78_N32574_O_4_C_2_io_in_WIRE_0 = IN_OPIN_N21942_38; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C78_N32574_O_4_C_2_io_in_lo = {IN_OPIN_N21958_54,IN_OPIN_N21950_46,IN_OPIN_N21942_38}; // @[TileFull.scala 207:13]
  wire  _SBMux_C78_N32574_O_4_C_2_io_in_WIRE_5 = IN_CHANX_N23556_96; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C78_N32574_O_4_C_2_io_in_WIRE_4 = IN_CHANX_N23446_78; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C78_N32574_O_4_C_2_io_in_hi_hi = {IN_CHANX_N23556_96,IN_CHANX_N23446_78}; // @[TileFull.scala 207:13]
  wire  _SBMux_C78_N32574_O_4_C_2_io_in_WIRE_3 = IN_OPIN_N21966_62; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C78_N32574_O_4_C_2_io_in_hi = {IN_CHANX_N23556_96,IN_CHANX_N23446_78,IN_OPIN_N21966_62}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C78_N32574_O_4_C_2_io_in_T = {IN_CHANX_N23556_96,IN_CHANX_N23446_78,IN_OPIN_N21966_62,
    IN_OPIN_N21958_54,IN_OPIN_N21950_46,IN_OPIN_N21942_38}; // @[TileFull.scala 207:13]
  wire  _SBMux_C80_N32576_O_4_C_2_io_in_WIRE_2 = IN_OPIN_N21959_55; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C80_N32576_O_4_C_2_io_in_WIRE_1 = IN_OPIN_N21951_47; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C80_N32576_O_4_C_2_io_in_lo_hi = {IN_OPIN_N21959_55,IN_OPIN_N21951_47}; // @[TileFull.scala 207:13]
  wire  _SBMux_C80_N32576_O_4_C_2_io_in_WIRE_0 = IN_OPIN_N21943_39; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C80_N32576_O_4_C_2_io_in_lo = {IN_OPIN_N21959_55,IN_OPIN_N21951_47,IN_OPIN_N21943_39}; // @[TileFull.scala 207:13]
  wire  _SBMux_C80_N32576_O_4_C_2_io_in_WIRE_5 = IN_CHANX_N23520_90; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C80_N32576_O_4_C_2_io_in_WIRE_4 = IN_CHANX_N23514_74; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C80_N32576_O_4_C_2_io_in_hi_hi = {IN_CHANX_N23520_90,IN_CHANX_N23514_74}; // @[TileFull.scala 207:13]
  wire  _SBMux_C80_N32576_O_4_C_2_io_in_WIRE_3 = IN_OPIN_N21967_63; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C80_N32576_O_4_C_2_io_in_hi = {IN_CHANX_N23520_90,IN_CHANX_N23514_74,IN_OPIN_N21967_63}; // @[TileFull.scala 207:13]
  wire [5:0] _SBMux_C80_N32576_O_4_C_2_io_in_T = {IN_CHANX_N23520_90,IN_CHANX_N23514_74,IN_OPIN_N21967_63,
    IN_OPIN_N21959_55,IN_OPIN_N21951_47,IN_OPIN_N21943_39}; // @[TileFull.scala 207:13]
  wire  _SBMux_C82_N32578_O_3_C_2_io_in_WIRE_1 = IN_OPIN_N21949_45; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C82_N32578_O_3_C_2_io_in_WIRE_0 = IN_OPIN_N21936_32; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C82_N32578_O_3_C_2_io_in_lo = {IN_OPIN_N21949_45,IN_OPIN_N21936_32}; // @[TileFull.scala 207:13]
  wire  _SBMux_C82_N32578_O_3_C_2_io_in_WIRE_4 = IN_CHANX_N23516_82; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C82_N32578_O_3_C_2_io_in_WIRE_3 = IN_CHANX_N23476_56; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C82_N32578_O_3_C_2_io_in_hi_hi = {IN_CHANX_N23516_82,IN_CHANX_N23476_56}; // @[TileFull.scala 207:13]
  wire  _SBMux_C82_N32578_O_3_C_2_io_in_WIRE_2 = IN_OPIN_N21962_58; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C82_N32578_O_3_C_2_io_in_hi = {IN_CHANX_N23516_82,IN_CHANX_N23476_56,IN_OPIN_N21962_58}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C82_N32578_O_3_C_2_io_in_T = {IN_CHANX_N23516_82,IN_CHANX_N23476_56,IN_OPIN_N21962_58,
    IN_OPIN_N21949_45,IN_OPIN_N21936_32}; // @[TileFull.scala 207:13]
  wire  _SBMux_C84_N32580_O_3_C_2_io_in_WIRE_1 = IN_OPIN_N21950_46; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C84_N32580_O_3_C_2_io_in_WIRE_0 = IN_OPIN_N21937_33; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C84_N32580_O_3_C_2_io_in_lo = {IN_OPIN_N21950_46,IN_OPIN_N21937_33}; // @[TileFull.scala 207:13]
  wire  _SBMux_C84_N32580_O_3_C_2_io_in_WIRE_4 = IN_CHANX_N23524_98; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C84_N32580_O_3_C_2_io_in_WIRE_3 = IN_CHANX_N23462_0; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C84_N32580_O_3_C_2_io_in_hi_hi = {IN_CHANX_N23524_98,IN_CHANX_N23462_0}; // @[TileFull.scala 207:13]
  wire  _SBMux_C84_N32580_O_3_C_2_io_in_WIRE_2 = IN_OPIN_N21963_59; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C84_N32580_O_3_C_2_io_in_hi = {IN_CHANX_N23524_98,IN_CHANX_N23462_0,IN_OPIN_N21963_59}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C84_N32580_O_3_C_2_io_in_T = {IN_CHANX_N23524_98,IN_CHANX_N23462_0,IN_OPIN_N21963_59,
    IN_OPIN_N21950_46,IN_OPIN_N21937_33}; // @[TileFull.scala 207:13]
  wire  _SBMux_C86_N32582_O_3_C_2_io_in_WIRE_1 = IN_OPIN_N21951_47; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C86_N32582_O_3_C_2_io_in_WIRE_0 = IN_OPIN_N21938_34; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C86_N32582_O_3_C_2_io_in_lo = {IN_OPIN_N21951_47,IN_OPIN_N21938_34}; // @[TileFull.scala 207:13]
  wire  _SBMux_C86_N32582_O_3_C_2_io_in_WIRE_4 = IN_CHANX_N23550_84; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C86_N32582_O_3_C_2_io_in_WIRE_3 = IN_CHANX_N23470_32; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C86_N32582_O_3_C_2_io_in_hi_hi = {IN_CHANX_N23550_84,IN_CHANX_N23470_32}; // @[TileFull.scala 207:13]
  wire  _SBMux_C86_N32582_O_3_C_2_io_in_WIRE_2 = IN_OPIN_N21964_60; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C86_N32582_O_3_C_2_io_in_hi = {IN_CHANX_N23550_84,IN_CHANX_N23470_32,IN_OPIN_N21964_60}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C86_N32582_O_3_C_2_io_in_T = {IN_CHANX_N23550_84,IN_CHANX_N23470_32,IN_OPIN_N21964_60,
    IN_OPIN_N21951_47,IN_OPIN_N21938_34}; // @[TileFull.scala 207:13]
  wire  _SBMux_C88_N32584_O_3_C_2_io_in_WIRE_1 = IN_OPIN_N21952_48; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C88_N32584_O_3_C_2_io_in_WIRE_0 = IN_OPIN_N21939_35; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C88_N32584_O_3_C_2_io_in_lo = {IN_OPIN_N21952_48,IN_OPIN_N21939_35}; // @[TileFull.scala 207:13]
  wire  _SBMux_C88_N32584_O_3_C_2_io_in_WIRE_4 = IN_CHANX_N23518_86; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C88_N32584_O_3_C_2_io_in_WIRE_3 = IN_CHANX_N23496_2; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C88_N32584_O_3_C_2_io_in_hi_hi = {IN_CHANX_N23518_86,IN_CHANX_N23496_2}; // @[TileFull.scala 207:13]
  wire  _SBMux_C88_N32584_O_3_C_2_io_in_WIRE_2 = IN_OPIN_N21965_61; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C88_N32584_O_3_C_2_io_in_hi = {IN_CHANX_N23518_86,IN_CHANX_N23496_2,IN_OPIN_N21965_61}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C88_N32584_O_3_C_2_io_in_T = {IN_CHANX_N23518_86,IN_CHANX_N23496_2,IN_OPIN_N21965_61,
    IN_OPIN_N21952_48,IN_OPIN_N21939_35}; // @[TileFull.scala 207:13]
  wire  _SBMux_C90_N32586_O_3_C_2_io_in_WIRE_1 = IN_OPIN_N21953_49; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C90_N32586_O_3_C_2_io_in_WIRE_0 = IN_OPIN_N21940_36; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C90_N32586_O_3_C_2_io_in_lo = {IN_OPIN_N21953_49,IN_OPIN_N21940_36}; // @[TileFull.scala 207:13]
  wire  _SBMux_C90_N32586_O_3_C_2_io_in_WIRE_4 = IN_CHANX_N23532_12; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C90_N32586_O_3_C_2_io_in_WIRE_3 = IN_CHANX_N23522_94; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C90_N32586_O_3_C_2_io_in_hi_hi = {IN_CHANX_N23532_12,IN_CHANX_N23522_94}; // @[TileFull.scala 207:13]
  wire  _SBMux_C90_N32586_O_3_C_2_io_in_WIRE_2 = IN_OPIN_N21966_62; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C90_N32586_O_3_C_2_io_in_hi = {IN_CHANX_N23532_12,IN_CHANX_N23522_94,IN_OPIN_N21966_62}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C90_N32586_O_3_C_2_io_in_T = {IN_CHANX_N23532_12,IN_CHANX_N23522_94,IN_OPIN_N21966_62,
    IN_OPIN_N21953_49,IN_OPIN_N21940_36}; // @[TileFull.scala 207:13]
  wire  _SBMux_C92_N32588_O_3_C_2_io_in_WIRE_1 = IN_OPIN_N21954_50; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C92_N32588_O_3_C_2_io_in_WIRE_0 = IN_OPIN_N21941_37; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C92_N32588_O_3_C_2_io_in_lo = {IN_OPIN_N21954_50,IN_OPIN_N21941_37}; // @[TileFull.scala 207:13]
  wire  _SBMux_C92_N32588_O_3_C_2_io_in_WIRE_4 = IN_CHANX_N23552_88; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C92_N32588_O_3_C_2_io_in_WIRE_3 = IN_CHANX_N23428_6; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C92_N32588_O_3_C_2_io_in_hi_hi = {IN_CHANX_N23552_88,IN_CHANX_N23428_6}; // @[TileFull.scala 207:13]
  wire  _SBMux_C92_N32588_O_3_C_2_io_in_WIRE_2 = IN_OPIN_N21967_63; // @[TileFull.scala 192:{39,39}]
  wire [2:0] SBMux_C92_N32588_O_3_C_2_io_in_hi = {IN_CHANX_N23552_88,IN_CHANX_N23428_6,IN_OPIN_N21967_63}; // @[TileFull.scala 207:13]
  wire [4:0] _SBMux_C92_N32588_O_3_C_2_io_in_T = {IN_CHANX_N23552_88,IN_CHANX_N23428_6,IN_OPIN_N21967_63,
    IN_OPIN_N21954_50,IN_OPIN_N21941_37}; // @[TileFull.scala 207:13]
  wire  _SBMux_C94_N32590_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21955_51; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C94_N32590_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21942_38; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C94_N32590_O_2_C_2_io_in_lo = {IN_OPIN_N21955_51,IN_OPIN_N21942_38}; // @[TileFull.scala 207:13]
  wire  _SBMux_C94_N32590_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23558_100; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C94_N32590_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23442_62; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C94_N32590_O_2_C_2_io_in_hi = {IN_CHANX_N23558_100,IN_CHANX_N23442_62}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C94_N32590_O_2_C_2_io_in_T = {IN_CHANX_N23558_100,IN_CHANX_N23442_62,IN_OPIN_N21955_51,
    IN_OPIN_N21942_38}; // @[TileFull.scala 207:13]
  wire  _SBMux_C96_N32592_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21956_52; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C96_N32592_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21943_39; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C96_N32592_O_2_C_2_io_in_lo = {IN_OPIN_N21956_52,IN_OPIN_N21943_39}; // @[TileFull.scala 207:13]
  wire  _SBMux_C96_N32592_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23560_104; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C96_N32592_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23500_18; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C96_N32592_O_2_C_2_io_in_hi = {IN_CHANX_N23560_104,IN_CHANX_N23500_18}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C96_N32592_O_2_C_2_io_in_T = {IN_CHANX_N23560_104,IN_CHANX_N23500_18,IN_OPIN_N21956_52,
    IN_OPIN_N21943_39}; // @[TileFull.scala 207:13]
  wire  _SBMux_C98_N32594_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21957_53; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C98_N32594_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21944_40; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C98_N32594_O_2_C_2_io_in_lo = {IN_OPIN_N21957_53,IN_OPIN_N21944_40}; // @[TileFull.scala 207:13]
  wire  _SBMux_C98_N32594_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23554_92; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C98_N32594_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23430_14; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C98_N32594_O_2_C_2_io_in_hi = {IN_CHANX_N23554_92,IN_CHANX_N23430_14}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C98_N32594_O_2_C_2_io_in_T = {IN_CHANX_N23554_92,IN_CHANX_N23430_14,IN_OPIN_N21957_53,
    IN_OPIN_N21944_40}; // @[TileFull.scala 207:13]
  wire  _SBMux_C100_N32596_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21958_54; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C100_N32596_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21945_41; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C100_N32596_O_2_C_2_io_in_lo = {IN_OPIN_N21958_54,IN_OPIN_N21945_41}; // @[TileFull.scala 207:13]
  wire  _SBMux_C100_N32596_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23528_106; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C100_N32596_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23432_22; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C100_N32596_O_2_C_2_io_in_hi = {IN_CHANX_N23528_106,IN_CHANX_N23432_22}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C100_N32596_O_2_C_2_io_in_T = {IN_CHANX_N23528_106,IN_CHANX_N23432_22,IN_OPIN_N21958_54,
    IN_OPIN_N21945_41}; // @[TileFull.scala 207:13]
  wire  _SBMux_C102_N32598_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21959_55; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C102_N32598_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21946_42; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C102_N32598_O_2_C_2_io_in_lo = {IN_OPIN_N21959_55,IN_OPIN_N21946_42}; // @[TileFull.scala 207:13]
  wire  _SBMux_C102_N32598_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23556_96; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C102_N32598_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23530_4; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C102_N32598_O_2_C_2_io_in_hi = {IN_CHANX_N23556_96,IN_CHANX_N23530_4}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C102_N32598_O_2_C_2_io_in_T = {IN_CHANX_N23556_96,IN_CHANX_N23530_4,IN_OPIN_N21959_55,
    IN_OPIN_N21946_42}; // @[TileFull.scala 207:13]
  wire  _SBMux_C104_N32600_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21960_56; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C104_N32600_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21947_43; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C104_N32600_O_2_C_2_io_in_lo = {IN_OPIN_N21960_56,IN_OPIN_N21947_43}; // @[TileFull.scala 207:13]
  wire  _SBMux_C104_N32600_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23520_90; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C104_N32600_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23478_64; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C104_N32600_O_2_C_2_io_in_hi = {IN_CHANX_N23520_90,IN_CHANX_N23478_64}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C104_N32600_O_2_C_2_io_in_T = {IN_CHANX_N23520_90,IN_CHANX_N23478_64,IN_OPIN_N21960_56,
    IN_OPIN_N21947_43}; // @[TileFull.scala 207:13]
  wire  _SBMux_C106_N32602_O_2_C_2_io_in_WIRE_1 = IN_OPIN_N21961_57; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C106_N32602_O_2_C_2_io_in_WIRE_0 = IN_OPIN_N21948_44; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C106_N32602_O_2_C_2_io_in_lo = {IN_OPIN_N21961_57,IN_OPIN_N21948_44}; // @[TileFull.scala 207:13]
  wire  _SBMux_C106_N32602_O_2_C_2_io_in_WIRE_3 = IN_CHANX_N23538_36; // @[TileFull.scala 192:{39,39}]
  wire  _SBMux_C106_N32602_O_2_C_2_io_in_WIRE_2 = IN_CHANX_N23526_102; // @[TileFull.scala 192:{39,39}]
  wire [1:0] SBMux_C106_N32602_O_2_C_2_io_in_hi = {IN_CHANX_N23538_36,IN_CHANX_N23526_102}; // @[TileFull.scala 207:13]
  wire [3:0] _SBMux_C106_N32602_O_2_C_2_io_in_T = {IN_CHANX_N23538_36,IN_CHANX_N23526_102,IN_OPIN_N21961_57,
    IN_OPIN_N21948_44}; // @[TileFull.scala 207:13]
  ScanConf_Tile_11_0_EMPTY configBlock ( // @[TileFull.scala 67:31]
    .clock(configBlock_clock),
    .reset(configBlock_reset),
    .ioBundle_confOut(configBlock_ioBundle_confOut),
    .ioBundle_scan_in(configBlock_ioBundle_scan_in),
    .ioBundle_scan_en(configBlock_ioBundle_scan_en),
    .ioBundle_scan_out(configBlock_ioBundle_scan_out),
    .ioBundle_scan_ioLatchEnb(configBlock_ioBundle_scan_ioLatchEnb)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C7_N23429_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C7_N23429_O_0_C_2_io_in),
    .io_config(SBMux_C7_N23429_O_0_C_2_io_config),
    .io_out(SBMux_C7_N23429_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C7_N23429_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C7_N23429_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C7_N23429_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C7_N23429_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C15_N23431_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C15_N23431_O_0_C_3_io_in),
    .io_config(SBMux_C15_N23431_O_0_C_3_io_config),
    .io_out(SBMux_C15_N23431_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C15_N23431_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C15_N23431_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C15_N23431_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C15_N23431_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C23_N23433_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C23_N23433_O_0_C_3_io_in),
    .io_config(SBMux_C23_N23433_O_0_C_3_io_config),
    .io_out(SBMux_C23_N23433_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C23_N23433_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C23_N23433_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C23_N23433_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C23_N23433_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C31_N23435_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C31_N23435_O_0_C_3_io_in),
    .io_config(SBMux_C31_N23435_O_0_C_3_io_config),
    .io_out(SBMux_C31_N23435_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C31_N23435_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C31_N23435_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C31_N23435_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C31_N23435_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C39_N23437_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C39_N23437_O_0_C_3_io_in),
    .io_config(SBMux_C39_N23437_O_0_C_3_io_config),
    .io_out(SBMux_C39_N23437_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C39_N23437_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C39_N23437_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C39_N23437_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C39_N23437_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C47_N23439_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C47_N23439_O_0_C_3_io_in),
    .io_config(SBMux_C47_N23439_O_0_C_3_io_config),
    .io_out(SBMux_C47_N23439_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C47_N23439_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C47_N23439_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C47_N23439_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C47_N23439_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C5_SCAOptSB SBMux_C55_N23441_O_0_C_5 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C55_N23441_O_0_C_5_io_in),
    .io_config(SBMux_C55_N23441_O_0_C_5_io_config),
    .io_out(SBMux_C55_N23441_O_0_C_5_io_out),
    .io_loopBreak(SBMux_C55_N23441_O_0_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C55_N23441_O_0_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C55_N23441_O_0_C_5_io_cnstClk),
    .io_arst(SBMux_C55_N23441_O_0_C_5_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C63_N23443_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C63_N23443_O_0_C_3_io_in),
    .io_config(SBMux_C63_N23443_O_0_C_3_io_config),
    .io_out(SBMux_C63_N23443_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C63_N23443_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C63_N23443_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C63_N23443_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C63_N23443_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C71_N23445_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C71_N23445_O_0_C_2_io_in),
    .io_config(SBMux_C71_N23445_O_0_C_2_io_config),
    .io_out(SBMux_C71_N23445_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C71_N23445_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C71_N23445_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C71_N23445_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C71_N23445_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C79_N23447_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C79_N23447_O_0_C_2_io_in),
    .io_config(SBMux_C79_N23447_O_0_C_2_io_config),
    .io_out(SBMux_C79_N23447_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C79_N23447_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C79_N23447_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C79_N23447_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C79_N23447_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C1_N23463_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C1_N23463_O_0_C_2_io_in),
    .io_config(SBMux_C1_N23463_O_0_C_2_io_config),
    .io_out(SBMux_C1_N23463_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C1_N23463_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C1_N23463_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C1_N23463_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C1_N23463_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C9_N23465_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C9_N23465_O_0_C_3_io_in),
    .io_config(SBMux_C9_N23465_O_0_C_3_io_config),
    .io_out(SBMux_C9_N23465_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C9_N23465_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C9_N23465_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C9_N23465_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C9_N23465_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C17_N23467_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C17_N23467_O_0_C_3_io_in),
    .io_config(SBMux_C17_N23467_O_0_C_3_io_config),
    .io_out(SBMux_C17_N23467_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C17_N23467_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C17_N23467_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C17_N23467_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C17_N23467_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C25_N23469_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C25_N23469_O_0_C_3_io_in),
    .io_config(SBMux_C25_N23469_O_0_C_3_io_config),
    .io_out(SBMux_C25_N23469_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C25_N23469_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C25_N23469_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C25_N23469_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C25_N23469_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C4_SCAOptSB SBMux_C33_N23471_O_0_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C33_N23471_O_0_C_4_io_in),
    .io_config(SBMux_C33_N23471_O_0_C_4_io_config),
    .io_out(SBMux_C33_N23471_O_0_C_4_io_out),
    .io_loopBreak(SBMux_C33_N23471_O_0_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C33_N23471_O_0_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C33_N23471_O_0_C_4_io_cnstClk),
    .io_arst(SBMux_C33_N23471_O_0_C_4_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C41_N23473_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C41_N23473_O_0_C_3_io_in),
    .io_config(SBMux_C41_N23473_O_0_C_3_io_config),
    .io_out(SBMux_C41_N23473_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C41_N23473_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C41_N23473_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C41_N23473_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C41_N23473_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C4_SCAOptSB SBMux_C49_N23475_O_0_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C49_N23475_O_0_C_4_io_in),
    .io_config(SBMux_C49_N23475_O_0_C_4_io_config),
    .io_out(SBMux_C49_N23475_O_0_C_4_io_out),
    .io_loopBreak(SBMux_C49_N23475_O_0_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C49_N23475_O_0_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C49_N23475_O_0_C_4_io_cnstClk),
    .io_arst(SBMux_C49_N23475_O_0_C_4_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C57_N23477_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C57_N23477_O_0_C_3_io_in),
    .io_config(SBMux_C57_N23477_O_0_C_3_io_config),
    .io_out(SBMux_C57_N23477_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C57_N23477_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C57_N23477_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C57_N23477_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C57_N23477_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C4_SCAOptSB SBMux_C65_N23479_O_0_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C65_N23479_O_0_C_4_io_in),
    .io_config(SBMux_C65_N23479_O_0_C_4_io_config),
    .io_out(SBMux_C65_N23479_O_0_C_4_io_out),
    .io_loopBreak(SBMux_C65_N23479_O_0_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C65_N23479_O_0_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C65_N23479_O_0_C_4_io_cnstClk),
    .io_arst(SBMux_C65_N23479_O_0_C_4_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C73_N23481_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C73_N23481_O_0_C_2_io_in),
    .io_config(SBMux_C73_N23481_O_0_C_2_io_config),
    .io_out(SBMux_C73_N23481_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C73_N23481_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C73_N23481_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C73_N23481_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C73_N23481_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C81_N23483_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C81_N23483_O_0_C_2_io_in),
    .io_config(SBMux_C81_N23483_O_0_C_2_io_config),
    .io_out(SBMux_C81_N23483_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C81_N23483_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C81_N23483_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C81_N23483_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C81_N23483_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C3_N23497_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C3_N23497_O_0_C_3_io_in),
    .io_config(SBMux_C3_N23497_O_0_C_3_io_config),
    .io_out(SBMux_C3_N23497_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C3_N23497_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C3_N23497_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C3_N23497_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C3_N23497_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C11_N23499_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C11_N23499_O_0_C_3_io_in),
    .io_config(SBMux_C11_N23499_O_0_C_3_io_config),
    .io_out(SBMux_C11_N23499_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C11_N23499_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C11_N23499_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C11_N23499_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C11_N23499_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C19_N23501_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C19_N23501_O_0_C_3_io_in),
    .io_config(SBMux_C19_N23501_O_0_C_3_io_config),
    .io_out(SBMux_C19_N23501_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C19_N23501_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C19_N23501_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C19_N23501_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C19_N23501_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C4_SCAOptSB SBMux_C27_N23503_O_0_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C27_N23503_O_0_C_4_io_in),
    .io_config(SBMux_C27_N23503_O_0_C_4_io_config),
    .io_out(SBMux_C27_N23503_O_0_C_4_io_out),
    .io_loopBreak(SBMux_C27_N23503_O_0_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C27_N23503_O_0_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C27_N23503_O_0_C_4_io_cnstClk),
    .io_arst(SBMux_C27_N23503_O_0_C_4_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C35_N23505_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C35_N23505_O_0_C_3_io_in),
    .io_config(SBMux_C35_N23505_O_0_C_3_io_config),
    .io_out(SBMux_C35_N23505_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C35_N23505_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C35_N23505_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C35_N23505_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C35_N23505_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C4_SCAOptSB SBMux_C43_N23507_O_0_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C43_N23507_O_0_C_4_io_in),
    .io_config(SBMux_C43_N23507_O_0_C_4_io_config),
    .io_out(SBMux_C43_N23507_O_0_C_4_io_out),
    .io_loopBreak(SBMux_C43_N23507_O_0_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C43_N23507_O_0_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C43_N23507_O_0_C_4_io_cnstClk),
    .io_arst(SBMux_C43_N23507_O_0_C_4_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C51_N23509_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C51_N23509_O_0_C_2_io_in),
    .io_config(SBMux_C51_N23509_O_0_C_2_io_config),
    .io_out(SBMux_C51_N23509_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C51_N23509_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C51_N23509_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C51_N23509_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C51_N23509_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C59_N23511_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C59_N23511_O_0_C_3_io_in),
    .io_config(SBMux_C59_N23511_O_0_C_3_io_config),
    .io_out(SBMux_C59_N23511_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C59_N23511_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C59_N23511_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C59_N23511_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C59_N23511_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C67_N23513_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C67_N23513_O_0_C_2_io_in),
    .io_config(SBMux_C67_N23513_O_0_C_2_io_config),
    .io_out(SBMux_C67_N23513_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C67_N23513_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C67_N23513_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C67_N23513_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C67_N23513_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C75_N23515_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C75_N23515_O_0_C_2_io_in),
    .io_config(SBMux_C75_N23515_O_0_C_2_io_config),
    .io_out(SBMux_C75_N23515_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C75_N23515_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C75_N23515_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C75_N23515_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C75_N23515_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C83_N23517_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C83_N23517_O_0_C_2_io_in),
    .io_config(SBMux_C83_N23517_O_0_C_2_io_config),
    .io_out(SBMux_C83_N23517_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C83_N23517_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C83_N23517_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C83_N23517_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C83_N23517_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C87_N23519_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C87_N23519_O_0_C_2_io_in),
    .io_config(SBMux_C87_N23519_O_0_C_2_io_config),
    .io_out(SBMux_C87_N23519_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C87_N23519_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C87_N23519_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C87_N23519_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C87_N23519_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C91_N23521_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C91_N23521_O_0_C_2_io_in),
    .io_config(SBMux_C91_N23521_O_0_C_2_io_config),
    .io_out(SBMux_C91_N23521_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C91_N23521_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C91_N23521_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C91_N23521_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C91_N23521_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C95_N23523_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C95_N23523_O_0_C_2_io_in),
    .io_config(SBMux_C95_N23523_O_0_C_2_io_config),
    .io_out(SBMux_C95_N23523_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C95_N23523_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C95_N23523_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C95_N23523_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C95_N23523_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C99_N23525_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C99_N23525_O_0_C_2_io_in),
    .io_config(SBMux_C99_N23525_O_0_C_2_io_config),
    .io_out(SBMux_C99_N23525_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C99_N23525_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C99_N23525_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C99_N23525_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C99_N23525_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C103_N23527_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C103_N23527_O_0_C_2_io_in),
    .io_config(SBMux_C103_N23527_O_0_C_2_io_config),
    .io_out(SBMux_C103_N23527_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C103_N23527_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C103_N23527_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C103_N23527_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C103_N23527_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C107_N23529_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C107_N23529_O_0_C_2_io_in),
    .io_config(SBMux_C107_N23529_O_0_C_2_io_config),
    .io_out(SBMux_C107_N23529_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C107_N23529_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C107_N23529_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C107_N23529_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C107_N23529_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C5_N23531_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C5_N23531_O_0_C_2_io_in),
    .io_config(SBMux_C5_N23531_O_0_C_2_io_config),
    .io_out(SBMux_C5_N23531_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C5_N23531_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C5_N23531_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C5_N23531_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C5_N23531_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C13_N23533_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C13_N23533_O_0_C_2_io_in),
    .io_config(SBMux_C13_N23533_O_0_C_2_io_config),
    .io_out(SBMux_C13_N23533_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C13_N23533_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C13_N23533_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C13_N23533_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C13_N23533_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C21_N23535_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C21_N23535_O_0_C_3_io_in),
    .io_config(SBMux_C21_N23535_O_0_C_3_io_config),
    .io_out(SBMux_C21_N23535_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C21_N23535_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C21_N23535_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C21_N23535_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C21_N23535_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C29_N23537_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C29_N23537_O_0_C_2_io_in),
    .io_config(SBMux_C29_N23537_O_0_C_2_io_config),
    .io_out(SBMux_C29_N23537_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C29_N23537_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C29_N23537_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C29_N23537_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C29_N23537_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C37_N23539_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C37_N23539_O_0_C_3_io_in),
    .io_config(SBMux_C37_N23539_O_0_C_3_io_config),
    .io_out(SBMux_C37_N23539_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C37_N23539_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C37_N23539_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C37_N23539_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C37_N23539_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C45_N23541_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C45_N23541_O_0_C_2_io_in),
    .io_config(SBMux_C45_N23541_O_0_C_2_io_config),
    .io_out(SBMux_C45_N23541_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C45_N23541_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C45_N23541_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C45_N23541_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C45_N23541_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C53_N23543_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C53_N23543_O_0_C_3_io_in),
    .io_config(SBMux_C53_N23543_O_0_C_3_io_config),
    .io_out(SBMux_C53_N23543_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C53_N23543_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C53_N23543_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C53_N23543_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C53_N23543_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C3_SCAOptSB SBMux_C61_N23545_O_0_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C61_N23545_O_0_C_3_io_in),
    .io_config(SBMux_C61_N23545_O_0_C_3_io_config),
    .io_out(SBMux_C61_N23545_O_0_C_3_io_out),
    .io_loopBreak(SBMux_C61_N23545_O_0_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C61_N23545_O_0_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C61_N23545_O_0_C_3_io_cnstClk),
    .io_arst(SBMux_C61_N23545_O_0_C_3_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C69_N23547_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C69_N23547_O_0_C_2_io_in),
    .io_config(SBMux_C69_N23547_O_0_C_2_io_config),
    .io_out(SBMux_C69_N23547_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C69_N23547_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C69_N23547_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C69_N23547_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C69_N23547_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C77_N23549_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C77_N23549_O_0_C_2_io_in),
    .io_config(SBMux_C77_N23549_O_0_C_2_io_config),
    .io_out(SBMux_C77_N23549_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C77_N23549_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C77_N23549_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C77_N23549_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C77_N23549_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C85_N23551_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C85_N23551_O_0_C_2_io_in),
    .io_config(SBMux_C85_N23551_O_0_C_2_io_config),
    .io_out(SBMux_C85_N23551_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C85_N23551_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C85_N23551_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C85_N23551_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C85_N23551_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C89_N23553_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C89_N23553_O_0_C_2_io_in),
    .io_config(SBMux_C89_N23553_O_0_C_2_io_config),
    .io_out(SBMux_C89_N23553_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C89_N23553_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C89_N23553_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C89_N23553_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C89_N23553_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C93_N23555_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C93_N23555_O_0_C_2_io_in),
    .io_config(SBMux_C93_N23555_O_0_C_2_io_config),
    .io_out(SBMux_C93_N23555_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C93_N23555_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C93_N23555_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C93_N23555_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C93_N23555_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C97_N23557_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C97_N23557_O_0_C_2_io_in),
    .io_config(SBMux_C97_N23557_O_0_C_2_io_config),
    .io_out(SBMux_C97_N23557_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C97_N23557_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C97_N23557_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C97_N23557_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C97_N23557_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C101_N23559_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C101_N23559_O_0_C_2_io_in),
    .io_config(SBMux_C101_N23559_O_0_C_2_io_config),
    .io_out(SBMux_C101_N23559_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C101_N23559_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C101_N23559_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C101_N23559_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C101_N23559_O_0_C_2_io_arst)
  );
  MuxNInput_O0_C2_SCAOptSB SBMux_C105_N23561_O_0_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C105_N23561_O_0_C_2_io_in),
    .io_config(SBMux_C105_N23561_O_0_C_2_io_config),
    .io_out(SBMux_C105_N23561_O_0_C_2_io_out),
    .io_loopBreak(SBMux_C105_N23561_O_0_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C105_N23561_O_0_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C105_N23561_O_0_C_2_io_cnstClk),
    .io_arst(SBMux_C105_N23561_O_0_C_2_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C0_N32496_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C0_N32496_O_2_C_3_io_in),
    .io_config(SBMux_C0_N32496_O_2_C_3_io_config),
    .io_out(SBMux_C0_N32496_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C0_N32496_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C0_N32496_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C0_N32496_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C0_N32496_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C2_N32498_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C2_N32498_O_2_C_3_io_in),
    .io_config(SBMux_C2_N32498_O_2_C_3_io_config),
    .io_out(SBMux_C2_N32498_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C2_N32498_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C2_N32498_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C2_N32498_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C2_N32498_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C4_N32500_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C4_N32500_O_2_C_3_io_in),
    .io_config(SBMux_C4_N32500_O_2_C_3_io_config),
    .io_out(SBMux_C4_N32500_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C4_N32500_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C4_N32500_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C4_N32500_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C4_N32500_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C4_SCAOptSB SBMux_C6_N32502_O_2_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C6_N32502_O_2_C_4_io_in),
    .io_config(SBMux_C6_N32502_O_2_C_4_io_config),
    .io_out(SBMux_C6_N32502_O_2_C_4_io_out),
    .io_loopBreak(SBMux_C6_N32502_O_2_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C6_N32502_O_2_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C6_N32502_O_2_C_4_io_cnstClk),
    .io_arst(SBMux_C6_N32502_O_2_C_4_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C8_N32504_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C8_N32504_O_2_C_3_io_in),
    .io_config(SBMux_C8_N32504_O_2_C_3_io_config),
    .io_out(SBMux_C8_N32504_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C8_N32504_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C8_N32504_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C8_N32504_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C8_N32504_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C4_SCAOptSB SBMux_C10_N32506_O_2_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C10_N32506_O_2_C_4_io_in),
    .io_config(SBMux_C10_N32506_O_2_C_4_io_config),
    .io_out(SBMux_C10_N32506_O_2_C_4_io_out),
    .io_loopBreak(SBMux_C10_N32506_O_2_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C10_N32506_O_2_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C10_N32506_O_2_C_4_io_cnstClk),
    .io_arst(SBMux_C10_N32506_O_2_C_4_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C12_N32508_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C12_N32508_O_2_C_3_io_in),
    .io_config(SBMux_C12_N32508_O_2_C_3_io_config),
    .io_out(SBMux_C12_N32508_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C12_N32508_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C12_N32508_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C12_N32508_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C12_N32508_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C4_SCAOptSB SBMux_C14_N32510_O_2_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C14_N32510_O_2_C_4_io_in),
    .io_config(SBMux_C14_N32510_O_2_C_4_io_config),
    .io_out(SBMux_C14_N32510_O_2_C_4_io_out),
    .io_loopBreak(SBMux_C14_N32510_O_2_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C14_N32510_O_2_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C14_N32510_O_2_C_4_io_cnstClk),
    .io_arst(SBMux_C14_N32510_O_2_C_4_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C16_N32512_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C16_N32512_O_2_C_3_io_in),
    .io_config(SBMux_C16_N32512_O_2_C_3_io_config),
    .io_out(SBMux_C16_N32512_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C16_N32512_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C16_N32512_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C16_N32512_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C16_N32512_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C4_SCAOptSB SBMux_C18_N32514_O_2_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C18_N32514_O_2_C_4_io_in),
    .io_config(SBMux_C18_N32514_O_2_C_4_io_config),
    .io_out(SBMux_C18_N32514_O_2_C_4_io_out),
    .io_loopBreak(SBMux_C18_N32514_O_2_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C18_N32514_O_2_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C18_N32514_O_2_C_4_io_cnstClk),
    .io_arst(SBMux_C18_N32514_O_2_C_4_io_arst)
  );
  MuxNInput_O2_C4_SCAOptSB SBMux_C20_N32516_O_2_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C20_N32516_O_2_C_4_io_in),
    .io_config(SBMux_C20_N32516_O_2_C_4_io_config),
    .io_out(SBMux_C20_N32516_O_2_C_4_io_out),
    .io_loopBreak(SBMux_C20_N32516_O_2_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C20_N32516_O_2_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C20_N32516_O_2_C_4_io_cnstClk),
    .io_arst(SBMux_C20_N32516_O_2_C_4_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C22_N32518_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C22_N32518_O_2_C_3_io_in),
    .io_config(SBMux_C22_N32518_O_2_C_3_io_config),
    .io_out(SBMux_C22_N32518_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C22_N32518_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C22_N32518_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C22_N32518_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C22_N32518_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C24_N32520_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C24_N32520_O_2_C_2_io_in),
    .io_config(SBMux_C24_N32520_O_2_C_2_io_config),
    .io_out(SBMux_C24_N32520_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C24_N32520_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C24_N32520_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C24_N32520_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C24_N32520_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C26_N32522_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C26_N32522_O_2_C_3_io_in),
    .io_config(SBMux_C26_N32522_O_2_C_3_io_config),
    .io_out(SBMux_C26_N32522_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C26_N32522_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C26_N32522_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C26_N32522_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C26_N32522_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C28_N32524_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C28_N32524_O_2_C_2_io_in),
    .io_config(SBMux_C28_N32524_O_2_C_2_io_config),
    .io_out(SBMux_C28_N32524_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C28_N32524_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C28_N32524_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C28_N32524_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C28_N32524_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C30_N32526_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C30_N32526_O_2_C_2_io_in),
    .io_config(SBMux_C30_N32526_O_2_C_2_io_config),
    .io_out(SBMux_C30_N32526_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C30_N32526_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C30_N32526_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C30_N32526_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C30_N32526_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C4_SCAOptSB SBMux_C32_N32528_O_2_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C32_N32528_O_2_C_4_io_in),
    .io_config(SBMux_C32_N32528_O_2_C_4_io_config),
    .io_out(SBMux_C32_N32528_O_2_C_4_io_out),
    .io_loopBreak(SBMux_C32_N32528_O_2_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C32_N32528_O_2_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C32_N32528_O_2_C_4_io_cnstClk),
    .io_arst(SBMux_C32_N32528_O_2_C_4_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C34_N32530_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C34_N32530_O_2_C_3_io_in),
    .io_config(SBMux_C34_N32530_O_2_C_3_io_config),
    .io_out(SBMux_C34_N32530_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C34_N32530_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C34_N32530_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C34_N32530_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C34_N32530_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C36_N32532_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C36_N32532_O_2_C_3_io_in),
    .io_config(SBMux_C36_N32532_O_2_C_3_io_config),
    .io_out(SBMux_C36_N32532_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C36_N32532_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C36_N32532_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C36_N32532_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C36_N32532_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C4_SCAOptSB SBMux_C38_N32534_O_2_C_4 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C38_N32534_O_2_C_4_io_in),
    .io_config(SBMux_C38_N32534_O_2_C_4_io_config),
    .io_out(SBMux_C38_N32534_O_2_C_4_io_out),
    .io_loopBreak(SBMux_C38_N32534_O_2_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C38_N32534_O_2_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C38_N32534_O_2_C_4_io_cnstClk),
    .io_arst(SBMux_C38_N32534_O_2_C_4_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C40_N32536_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C40_N32536_O_2_C_2_io_in),
    .io_config(SBMux_C40_N32536_O_2_C_2_io_config),
    .io_out(SBMux_C40_N32536_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C40_N32536_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C40_N32536_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C40_N32536_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C40_N32536_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C42_N32538_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C42_N32538_O_2_C_3_io_in),
    .io_config(SBMux_C42_N32538_O_2_C_3_io_config),
    .io_out(SBMux_C42_N32538_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C42_N32538_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C42_N32538_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C42_N32538_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C42_N32538_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C44_N32540_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C44_N32540_O_2_C_3_io_in),
    .io_config(SBMux_C44_N32540_O_2_C_3_io_config),
    .io_out(SBMux_C44_N32540_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C44_N32540_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C44_N32540_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C44_N32540_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C44_N32540_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C46_N32542_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C46_N32542_O_2_C_3_io_in),
    .io_config(SBMux_C46_N32542_O_2_C_3_io_config),
    .io_out(SBMux_C46_N32542_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C46_N32542_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C46_N32542_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C46_N32542_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C46_N32542_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C48_N32544_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C48_N32544_O_2_C_3_io_in),
    .io_config(SBMux_C48_N32544_O_2_C_3_io_config),
    .io_out(SBMux_C48_N32544_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C48_N32544_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C48_N32544_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C48_N32544_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C48_N32544_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C50_N32546_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C50_N32546_O_2_C_3_io_in),
    .io_config(SBMux_C50_N32546_O_2_C_3_io_config),
    .io_out(SBMux_C50_N32546_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C50_N32546_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C50_N32546_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C50_N32546_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C50_N32546_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C52_N32548_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C52_N32548_O_2_C_3_io_in),
    .io_config(SBMux_C52_N32548_O_2_C_3_io_config),
    .io_out(SBMux_C52_N32548_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C52_N32548_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C52_N32548_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C52_N32548_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C52_N32548_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C54_N32550_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C54_N32550_O_2_C_2_io_in),
    .io_config(SBMux_C54_N32550_O_2_C_2_io_config),
    .io_out(SBMux_C54_N32550_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C54_N32550_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C54_N32550_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C54_N32550_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C54_N32550_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C56_N32552_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C56_N32552_O_2_C_3_io_in),
    .io_config(SBMux_C56_N32552_O_2_C_3_io_config),
    .io_out(SBMux_C56_N32552_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C56_N32552_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C56_N32552_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C56_N32552_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C56_N32552_O_2_C_3_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C58_N32554_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C58_N32554_O_2_C_2_io_in),
    .io_config(SBMux_C58_N32554_O_2_C_2_io_config),
    .io_out(SBMux_C58_N32554_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C58_N32554_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C58_N32554_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C58_N32554_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C58_N32554_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C3_SCAOptSB SBMux_C60_N32556_O_2_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C60_N32556_O_2_C_3_io_in),
    .io_config(SBMux_C60_N32556_O_2_C_3_io_config),
    .io_out(SBMux_C60_N32556_O_2_C_3_io_out),
    .io_loopBreak(SBMux_C60_N32556_O_2_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C60_N32556_O_2_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C60_N32556_O_2_C_3_io_cnstClk),
    .io_arst(SBMux_C60_N32556_O_2_C_3_io_arst)
  );
  MuxNInput_O1_C3_SCAOptSB SBMux_C62_N32558_O_1_C_3 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C62_N32558_O_1_C_3_io_in),
    .io_config(SBMux_C62_N32558_O_1_C_3_io_config),
    .io_out(SBMux_C62_N32558_O_1_C_3_io_out),
    .io_loopBreak(SBMux_C62_N32558_O_1_C_3_io_loopBreak),
    .io_ioGndBle(SBMux_C62_N32558_O_1_C_3_io_ioGndBle),
    .io_cnstClk(SBMux_C62_N32558_O_1_C_3_io_cnstClk),
    .io_arst(SBMux_C62_N32558_O_1_C_3_io_arst)
  );
  MuxNInput_O1_C2_SCAOptSB SBMux_C64_N32560_O_1_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C64_N32560_O_1_C_2_io_in),
    .io_config(SBMux_C64_N32560_O_1_C_2_io_config),
    .io_out(SBMux_C64_N32560_O_1_C_2_io_out),
    .io_loopBreak(SBMux_C64_N32560_O_1_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C64_N32560_O_1_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C64_N32560_O_1_C_2_io_cnstClk),
    .io_arst(SBMux_C64_N32560_O_1_C_2_io_arst)
  );
  MuxNInput_O4_C2_SCAOptSB SBMux_C66_N32562_O_4_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C66_N32562_O_4_C_2_io_in),
    .io_config(SBMux_C66_N32562_O_4_C_2_io_config),
    .io_out(SBMux_C66_N32562_O_4_C_2_io_out),
    .io_loopBreak(SBMux_C66_N32562_O_4_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C66_N32562_O_4_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C66_N32562_O_4_C_2_io_cnstClk),
    .io_arst(SBMux_C66_N32562_O_4_C_2_io_arst)
  );
  MuxNInput_O4_C2_SCAOptSB SBMux_C68_N32564_O_4_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C68_N32564_O_4_C_2_io_in),
    .io_config(SBMux_C68_N32564_O_4_C_2_io_config),
    .io_out(SBMux_C68_N32564_O_4_C_2_io_out),
    .io_loopBreak(SBMux_C68_N32564_O_4_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C68_N32564_O_4_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C68_N32564_O_4_C_2_io_cnstClk),
    .io_arst(SBMux_C68_N32564_O_4_C_2_io_arst)
  );
  MuxNInput_O4_C2_SCAOptSB SBMux_C70_N32566_O_4_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C70_N32566_O_4_C_2_io_in),
    .io_config(SBMux_C70_N32566_O_4_C_2_io_config),
    .io_out(SBMux_C70_N32566_O_4_C_2_io_out),
    .io_loopBreak(SBMux_C70_N32566_O_4_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C70_N32566_O_4_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C70_N32566_O_4_C_2_io_cnstClk),
    .io_arst(SBMux_C70_N32566_O_4_C_2_io_arst)
  );
  MuxNInput_O4_C2_SCAOptSB SBMux_C72_N32568_O_4_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C72_N32568_O_4_C_2_io_in),
    .io_config(SBMux_C72_N32568_O_4_C_2_io_config),
    .io_out(SBMux_C72_N32568_O_4_C_2_io_out),
    .io_loopBreak(SBMux_C72_N32568_O_4_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C72_N32568_O_4_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C72_N32568_O_4_C_2_io_cnstClk),
    .io_arst(SBMux_C72_N32568_O_4_C_2_io_arst)
  );
  MuxNInput_O4_C2_SCAOptSB SBMux_C74_N32570_O_4_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C74_N32570_O_4_C_2_io_in),
    .io_config(SBMux_C74_N32570_O_4_C_2_io_config),
    .io_out(SBMux_C74_N32570_O_4_C_2_io_out),
    .io_loopBreak(SBMux_C74_N32570_O_4_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C74_N32570_O_4_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C74_N32570_O_4_C_2_io_cnstClk),
    .io_arst(SBMux_C74_N32570_O_4_C_2_io_arst)
  );
  MuxNInput_O4_C2_SCAOptSB SBMux_C76_N32572_O_4_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C76_N32572_O_4_C_2_io_in),
    .io_config(SBMux_C76_N32572_O_4_C_2_io_config),
    .io_out(SBMux_C76_N32572_O_4_C_2_io_out),
    .io_loopBreak(SBMux_C76_N32572_O_4_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C76_N32572_O_4_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C76_N32572_O_4_C_2_io_cnstClk),
    .io_arst(SBMux_C76_N32572_O_4_C_2_io_arst)
  );
  MuxNInput_O4_C2_SCAOptSB SBMux_C78_N32574_O_4_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C78_N32574_O_4_C_2_io_in),
    .io_config(SBMux_C78_N32574_O_4_C_2_io_config),
    .io_out(SBMux_C78_N32574_O_4_C_2_io_out),
    .io_loopBreak(SBMux_C78_N32574_O_4_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C78_N32574_O_4_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C78_N32574_O_4_C_2_io_cnstClk),
    .io_arst(SBMux_C78_N32574_O_4_C_2_io_arst)
  );
  MuxNInput_O4_C2_SCAOptSB SBMux_C80_N32576_O_4_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C80_N32576_O_4_C_2_io_in),
    .io_config(SBMux_C80_N32576_O_4_C_2_io_config),
    .io_out(SBMux_C80_N32576_O_4_C_2_io_out),
    .io_loopBreak(SBMux_C80_N32576_O_4_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C80_N32576_O_4_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C80_N32576_O_4_C_2_io_cnstClk),
    .io_arst(SBMux_C80_N32576_O_4_C_2_io_arst)
  );
  MuxNInput_O3_C2_SCAOptSB SBMux_C82_N32578_O_3_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C82_N32578_O_3_C_2_io_in),
    .io_config(SBMux_C82_N32578_O_3_C_2_io_config),
    .io_out(SBMux_C82_N32578_O_3_C_2_io_out),
    .io_loopBreak(SBMux_C82_N32578_O_3_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C82_N32578_O_3_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C82_N32578_O_3_C_2_io_cnstClk),
    .io_arst(SBMux_C82_N32578_O_3_C_2_io_arst)
  );
  MuxNInput_O3_C2_SCAOptSB SBMux_C84_N32580_O_3_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C84_N32580_O_3_C_2_io_in),
    .io_config(SBMux_C84_N32580_O_3_C_2_io_config),
    .io_out(SBMux_C84_N32580_O_3_C_2_io_out),
    .io_loopBreak(SBMux_C84_N32580_O_3_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C84_N32580_O_3_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C84_N32580_O_3_C_2_io_cnstClk),
    .io_arst(SBMux_C84_N32580_O_3_C_2_io_arst)
  );
  MuxNInput_O3_C2_SCAOptSB SBMux_C86_N32582_O_3_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C86_N32582_O_3_C_2_io_in),
    .io_config(SBMux_C86_N32582_O_3_C_2_io_config),
    .io_out(SBMux_C86_N32582_O_3_C_2_io_out),
    .io_loopBreak(SBMux_C86_N32582_O_3_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C86_N32582_O_3_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C86_N32582_O_3_C_2_io_cnstClk),
    .io_arst(SBMux_C86_N32582_O_3_C_2_io_arst)
  );
  MuxNInput_O3_C2_SCAOptSB SBMux_C88_N32584_O_3_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C88_N32584_O_3_C_2_io_in),
    .io_config(SBMux_C88_N32584_O_3_C_2_io_config),
    .io_out(SBMux_C88_N32584_O_3_C_2_io_out),
    .io_loopBreak(SBMux_C88_N32584_O_3_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C88_N32584_O_3_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C88_N32584_O_3_C_2_io_cnstClk),
    .io_arst(SBMux_C88_N32584_O_3_C_2_io_arst)
  );
  MuxNInput_O3_C2_SCAOptSB SBMux_C90_N32586_O_3_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C90_N32586_O_3_C_2_io_in),
    .io_config(SBMux_C90_N32586_O_3_C_2_io_config),
    .io_out(SBMux_C90_N32586_O_3_C_2_io_out),
    .io_loopBreak(SBMux_C90_N32586_O_3_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C90_N32586_O_3_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C90_N32586_O_3_C_2_io_cnstClk),
    .io_arst(SBMux_C90_N32586_O_3_C_2_io_arst)
  );
  MuxNInput_O3_C2_SCAOptSB SBMux_C92_N32588_O_3_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C92_N32588_O_3_C_2_io_in),
    .io_config(SBMux_C92_N32588_O_3_C_2_io_config),
    .io_out(SBMux_C92_N32588_O_3_C_2_io_out),
    .io_loopBreak(SBMux_C92_N32588_O_3_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C92_N32588_O_3_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C92_N32588_O_3_C_2_io_cnstClk),
    .io_arst(SBMux_C92_N32588_O_3_C_2_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C94_N32590_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C94_N32590_O_2_C_2_io_in),
    .io_config(SBMux_C94_N32590_O_2_C_2_io_config),
    .io_out(SBMux_C94_N32590_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C94_N32590_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C94_N32590_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C94_N32590_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C94_N32590_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C96_N32592_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C96_N32592_O_2_C_2_io_in),
    .io_config(SBMux_C96_N32592_O_2_C_2_io_config),
    .io_out(SBMux_C96_N32592_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C96_N32592_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C96_N32592_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C96_N32592_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C96_N32592_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C98_N32594_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C98_N32594_O_2_C_2_io_in),
    .io_config(SBMux_C98_N32594_O_2_C_2_io_config),
    .io_out(SBMux_C98_N32594_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C98_N32594_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C98_N32594_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C98_N32594_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C98_N32594_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C100_N32596_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C100_N32596_O_2_C_2_io_in),
    .io_config(SBMux_C100_N32596_O_2_C_2_io_config),
    .io_out(SBMux_C100_N32596_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C100_N32596_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C100_N32596_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C100_N32596_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C100_N32596_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C102_N32598_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C102_N32598_O_2_C_2_io_in),
    .io_config(SBMux_C102_N32598_O_2_C_2_io_config),
    .io_out(SBMux_C102_N32598_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C102_N32598_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C102_N32598_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C102_N32598_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C102_N32598_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C104_N32600_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C104_N32600_O_2_C_2_io_in),
    .io_config(SBMux_C104_N32600_O_2_C_2_io_config),
    .io_out(SBMux_C104_N32600_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C104_N32600_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C104_N32600_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C104_N32600_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C104_N32600_O_2_C_2_io_arst)
  );
  MuxNInput_O2_C2_SCAOptSB SBMux_C106_N32602_O_2_C_2 ( // @[TileFull.scala 146:27]
    .io_in(SBMux_C106_N32602_O_2_C_2_io_in),
    .io_config(SBMux_C106_N32602_O_2_C_2_io_config),
    .io_out(SBMux_C106_N32602_O_2_C_2_io_out),
    .io_loopBreak(SBMux_C106_N32602_O_2_C_2_io_loopBreak),
    .io_ioGndBle(SBMux_C106_N32602_O_2_C_2_io_ioGndBle),
    .io_cnstClk(SBMux_C106_N32602_O_2_C_2_io_cnstClk),
    .io_arst(SBMux_C106_N32602_O_2_C_2_io_arst)
  );
  assign OUT_CHANY_N32528_32 = SBMux_C32_N32528_O_2_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32584_88 = SBMux_C88_N32584_O_3_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32566_70 = SBMux_C70_N32566_O_4_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23429_7 = SBMux_C7_N23429_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23537_29 = SBMux_C29_N23537_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23553_89 = SBMux_C89_N23553_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32568_72 = SBMux_C72_N32568_O_4_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23523_95 = SBMux_C95_N23523_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32534_38 = SBMux_C38_N32534_O_2_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32586_90 = SBMux_C90_N32586_O_3_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32546_50 = SBMux_C50_N32546_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32512_16 = SBMux_C16_N32512_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32554_58 = SBMux_C58_N32554_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23505_35 = SBMux_C35_N23505_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32548_52 = SBMux_C52_N32548_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23543_53 = SBMux_C53_N23543_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32596_100 = SBMux_C100_N32596_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32594_98 = SBMux_C98_N32594_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32560_64 = SBMux_C64_N32560_O_1_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23521_91 = SBMux_C91_N23521_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32582_86 = SBMux_C86_N32582_O_3_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32598_102 = SBMux_C102_N32598_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23527_103 = SBMux_C103_N23527_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23551_85 = SBMux_C85_N23551_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32508_12 = SBMux_C12_N32508_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32570_74 = SBMux_C74_N32570_O_4_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23499_11 = SBMux_C11_N23499_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32502_6 = SBMux_C6_N32502_O_2_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23535_21 = SBMux_C21_N23535_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23525_99 = SBMux_C99_N23525_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23501_19 = SBMux_C19_N23501_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32580_84 = SBMux_C84_N32580_O_3_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23517_83 = SBMux_C83_N23517_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23531_5 = SBMux_C5_N23531_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32524_28 = SBMux_C28_N32524_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32532_36 = SBMux_C36_N32532_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32602_106 = SBMux_C106_N32602_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23477_57 = SBMux_C57_N23477_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23473_41 = SBMux_C41_N23473_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23479_65 = SBMux_C65_N23479_O_0_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32552_56 = SBMux_C56_N32552_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23555_93 = SBMux_C93_N23555_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23447_79 = SBMux_C79_N23447_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32592_96 = SBMux_C96_N32592_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23561_105 = SBMux_C105_N23561_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32522_26 = SBMux_C26_N32522_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23513_67 = SBMux_C67_N23513_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32510_14 = SBMux_C14_N32510_O_2_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32544_48 = SBMux_C48_N32544_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23431_15 = SBMux_C15_N23431_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23435_31 = SBMux_C31_N23435_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23503_27 = SBMux_C27_N23503_O_0_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32518_22 = SBMux_C22_N32518_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23463_1 = SBMux_C1_N23463_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23437_39 = SBMux_C39_N23437_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32530_34 = SBMux_C34_N32530_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32496_0 = SBMux_C0_N32496_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23529_107 = SBMux_C107_N23529_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23469_25 = SBMux_C25_N23469_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32588_92 = SBMux_C92_N32588_O_3_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32536_40 = SBMux_C40_N32536_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32574_78 = SBMux_C78_N32574_O_4_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32578_82 = SBMux_C82_N32578_O_3_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23475_49 = SBMux_C49_N23475_O_0_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32550_54 = SBMux_C54_N32550_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23443_63 = SBMux_C63_N23443_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32564_68 = SBMux_C68_N32564_O_4_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23467_17 = SBMux_C17_N23467_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23471_33 = SBMux_C33_N23471_O_0_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23433_23 = SBMux_C23_N23433_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32558_62 = SBMux_C62_N32558_O_1_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23559_101 = SBMux_C101_N23559_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32516_20 = SBMux_C20_N32516_O_2_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23549_77 = SBMux_C77_N23549_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32526_30 = SBMux_C30_N32526_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32500_4 = SBMux_C4_N32500_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23445_71 = SBMux_C71_N23445_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32498_2 = SBMux_C2_N32498_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23481_73 = SBMux_C73_N23481_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32540_44 = SBMux_C44_N32540_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23539_37 = SBMux_C37_N23539_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32506_10 = SBMux_C10_N32506_O_2_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23465_9 = SBMux_C9_N23465_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23483_81 = SBMux_C81_N23483_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23439_47 = SBMux_C47_N23439_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32576_80 = SBMux_C80_N32576_O_4_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23545_61 = SBMux_C61_N23545_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23515_75 = SBMux_C75_N23515_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32520_24 = SBMux_C24_N32520_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23497_3 = SBMux_C3_N23497_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23509_51 = SBMux_C51_N23509_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23541_45 = SBMux_C45_N23541_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32538_42 = SBMux_C42_N32538_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32542_46 = SBMux_C46_N32542_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32572_76 = SBMux_C76_N32572_O_4_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23507_43 = SBMux_C43_N23507_O_0_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32504_8 = SBMux_C8_N32504_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32600_104 = SBMux_C104_N32600_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32556_60 = SBMux_C60_N32556_O_2_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32590_94 = SBMux_C94_N32590_O_2_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32514_18 = SBMux_C18_N32514_O_2_C_4_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANY_N32562_66 = SBMux_C66_N32562_O_4_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23511_59 = SBMux_C59_N23511_O_0_C_3_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23441_55 = SBMux_C55_N23441_O_0_C_5_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23519_87 = SBMux_C87_N23519_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23533_13 = SBMux_C13_N23533_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23557_97 = SBMux_C97_N23557_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign OUT_CHANX_N23547_69 = SBMux_C69_N23547_O_0_C_2_io_out; // @[TileFull.scala 151:25]
  assign ioConf_confOut = configBlock_ioBundle_confOut[282:0]; // @[TileFull.scala 78:12]
  assign ioConf_scan_out = configBlock_ioBundle_scan_out; // @[TileFull.scala 78:12]
  assign configBlock_clock = ctrlSignals_confClock; // @[TileFull.scala 79:27]
  assign configBlock_reset = reset;
  assign configBlock_ioBundle_scan_in = ioConf_scan_in; // @[TileFull.scala 78:12]
  assign configBlock_ioBundle_scan_en = ioConf_scan_en; // @[TileFull.scala 78:12]
  assign configBlock_ioBundle_scan_ioLatchEnb = ioConf_scan_ioLatchEnb; // @[TileFull.scala 78:12]
  assign SBMux_C7_N23429_O_0_C_2_io_in = {IN_CHANY_N32569_73,IN_CHANY_N32529_33}; // @[TileFull.scala 207:13]
  assign SBMux_C7_N23429_O_0_C_2_io_config = configBlock_ioBundle_confOut[1:0]; // @[TileFull.scala 156:60]
  assign SBMux_C7_N23429_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C7_N23429_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C7_N23429_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C7_N23429_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C15_N23431_O_0_C_3_io_in = {SBMux_C15_N23431_O_0_C_3_io_in_hi,IN_CHANY_N32509_13}; // @[TileFull.scala 207:13]
  assign SBMux_C15_N23431_O_0_C_3_io_config = configBlock_ioBundle_confOut[4:2]; // @[TileFull.scala 156:60]
  assign SBMux_C15_N23431_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C15_N23431_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C15_N23431_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C15_N23431_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C23_N23433_O_0_C_3_io_in = {SBMux_C23_N23433_O_0_C_3_io_in_hi,IN_CHANY_N32505_9}; // @[TileFull.scala 207:13]
  assign SBMux_C23_N23433_O_0_C_3_io_config = configBlock_ioBundle_confOut[7:5]; // @[TileFull.scala 156:60]
  assign SBMux_C23_N23433_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C23_N23433_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C23_N23433_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C23_N23433_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C31_N23435_O_0_C_3_io_in = {SBMux_C31_N23435_O_0_C_3_io_in_hi,IN_CHANY_N32561_65}; // @[TileFull.scala 207:13]
  assign SBMux_C31_N23435_O_0_C_3_io_config = configBlock_ioBundle_confOut[10:8]; // @[TileFull.scala 156:60]
  assign SBMux_C31_N23435_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C31_N23435_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C31_N23435_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C31_N23435_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C39_N23437_O_0_C_3_io_in = {SBMux_C39_N23437_O_0_C_3_io_in_hi,IN_CHANY_N32513_17}; // @[TileFull.scala 207:13]
  assign SBMux_C39_N23437_O_0_C_3_io_config = configBlock_ioBundle_confOut[13:11]; // @[TileFull.scala 156:60]
  assign SBMux_C39_N23437_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C39_N23437_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C39_N23437_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C39_N23437_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C47_N23439_O_0_C_3_io_in = {SBMux_C47_N23439_O_0_C_3_io_in_hi,IN_CHANY_N32535_39}; // @[TileFull.scala 207:13]
  assign SBMux_C47_N23439_O_0_C_3_io_config = configBlock_ioBundle_confOut[16:14]; // @[TileFull.scala 156:60]
  assign SBMux_C47_N23439_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C47_N23439_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C47_N23439_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C47_N23439_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C55_N23441_O_0_C_5_io_in = {SBMux_C55_N23441_O_0_C_5_io_in_hi,SBMux_C55_N23441_O_0_C_5_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C55_N23441_O_0_C_5_io_config = configBlock_ioBundle_confOut[20:17]; // @[TileFull.scala 156:60]
  assign SBMux_C55_N23441_O_0_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C55_N23441_O_0_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C55_N23441_O_0_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C55_N23441_O_0_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C63_N23443_O_0_C_3_io_in = {SBMux_C63_N23443_O_0_C_3_io_in_hi,IN_CHANY_N32511_15}; // @[TileFull.scala 207:13]
  assign SBMux_C63_N23443_O_0_C_3_io_config = configBlock_ioBundle_confOut[23:21]; // @[TileFull.scala 156:60]
  assign SBMux_C63_N23443_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C63_N23443_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C63_N23443_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C63_N23443_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C71_N23445_O_0_C_2_io_in = {IN_CHANY_N32599_103,IN_CHANY_N32567_71}; // @[TileFull.scala 207:13]
  assign SBMux_C71_N23445_O_0_C_2_io_config = configBlock_ioBundle_confOut[25:24]; // @[TileFull.scala 156:60]
  assign SBMux_C71_N23445_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C71_N23445_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C71_N23445_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C71_N23445_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C79_N23447_O_0_C_2_io_in = {IN_CHANY_N32597_101,IN_CHANY_N32563_67}; // @[TileFull.scala 207:13]
  assign SBMux_C79_N23447_O_0_C_2_io_config = configBlock_ioBundle_confOut[27:26]; // @[TileFull.scala 156:60]
  assign SBMux_C79_N23447_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C79_N23447_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C79_N23447_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C79_N23447_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C1_N23463_O_0_C_2_io_in = {IN_CHANY_N32575_79,IN_CHANY_N32531_35}; // @[TileFull.scala 207:13]
  assign SBMux_C1_N23463_O_0_C_2_io_config = configBlock_ioBundle_confOut[29:28]; // @[TileFull.scala 156:60]
  assign SBMux_C1_N23463_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C1_N23463_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C1_N23463_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C1_N23463_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C9_N23465_O_0_C_3_io_in = {SBMux_C9_N23465_O_0_C_3_io_in_hi,IN_CHANY_N32501_5}; // @[TileFull.scala 207:13]
  assign SBMux_C9_N23465_O_0_C_3_io_config = configBlock_ioBundle_confOut[32:30]; // @[TileFull.scala 156:60]
  assign SBMux_C9_N23465_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C9_N23465_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C9_N23465_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C9_N23465_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C17_N23467_O_0_C_3_io_in = {SBMux_C17_N23467_O_0_C_3_io_in_hi,IN_CHANY_N32559_63}; // @[TileFull.scala 207:13]
  assign SBMux_C17_N23467_O_0_C_3_io_config = configBlock_ioBundle_confOut[35:33]; // @[TileFull.scala 156:60]
  assign SBMux_C17_N23467_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C17_N23467_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C17_N23467_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C17_N23467_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C25_N23469_O_0_C_3_io_in = {SBMux_C25_N23469_O_0_C_3_io_in_hi,IN_CHANY_N32555_59}; // @[TileFull.scala 207:13]
  assign SBMux_C25_N23469_O_0_C_3_io_config = configBlock_ioBundle_confOut[38:36]; // @[TileFull.scala 156:60]
  assign SBMux_C25_N23469_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C25_N23469_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C25_N23469_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C25_N23469_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C33_N23471_O_0_C_4_io_in = {SBMux_C33_N23471_O_0_C_4_io_in_hi,SBMux_C33_N23471_O_0_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C33_N23471_O_0_C_4_io_config = configBlock_ioBundle_confOut[41:39]; // @[TileFull.scala 156:60]
  assign SBMux_C33_N23471_O_0_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C33_N23471_O_0_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C33_N23471_O_0_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C33_N23471_O_0_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C41_N23473_O_0_C_3_io_in = {SBMux_C41_N23473_O_0_C_3_io_in_hi,IN_CHANY_N32541_45}; // @[TileFull.scala 207:13]
  assign SBMux_C41_N23473_O_0_C_3_io_config = configBlock_ioBundle_confOut[44:42]; // @[TileFull.scala 156:60]
  assign SBMux_C41_N23473_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C41_N23473_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C41_N23473_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C41_N23473_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C49_N23475_O_0_C_4_io_in = {SBMux_C49_N23475_O_0_C_4_io_in_hi,SBMux_C49_N23475_O_0_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C49_N23475_O_0_C_4_io_config = configBlock_ioBundle_confOut[47:45]; // @[TileFull.scala 156:60]
  assign SBMux_C49_N23475_O_0_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C49_N23475_O_0_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C49_N23475_O_0_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C49_N23475_O_0_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C57_N23477_O_0_C_3_io_in = {SBMux_C57_N23477_O_0_C_3_io_in_hi,IN_CHANY_N32499_3}; // @[TileFull.scala 207:13]
  assign SBMux_C57_N23477_O_0_C_3_io_config = configBlock_ioBundle_confOut[50:48]; // @[TileFull.scala 156:60]
  assign SBMux_C57_N23477_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C57_N23477_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C57_N23477_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C57_N23477_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C65_N23479_O_0_C_4_io_in = {SBMux_C65_N23479_O_0_C_4_io_in_hi,SBMux_C65_N23479_O_0_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C65_N23479_O_0_C_4_io_config = configBlock_ioBundle_confOut[53:51]; // @[TileFull.scala 156:60]
  assign SBMux_C65_N23479_O_0_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C65_N23479_O_0_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C65_N23479_O_0_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C65_N23479_O_0_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C73_N23481_O_0_C_2_io_in = {IN_CHANY_N32585_89,IN_CHANY_N32565_69}; // @[TileFull.scala 207:13]
  assign SBMux_C73_N23481_O_0_C_2_io_config = configBlock_ioBundle_confOut[55:54]; // @[TileFull.scala 156:60]
  assign SBMux_C73_N23481_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C73_N23481_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C73_N23481_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C73_N23481_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C81_N23483_O_0_C_2_io_in = {IN_CHANY_N32595_99,IN_CHANY_N32577_81}; // @[TileFull.scala 207:13]
  assign SBMux_C81_N23483_O_0_C_2_io_config = configBlock_ioBundle_confOut[57:56]; // @[TileFull.scala 156:60]
  assign SBMux_C81_N23483_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C81_N23483_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C81_N23483_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C81_N23483_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C3_N23497_O_0_C_3_io_in = {SBMux_C3_N23497_O_0_C_3_io_in_hi,IN_CHANY_N32525_29}; // @[TileFull.scala 207:13]
  assign SBMux_C3_N23497_O_0_C_3_io_config = configBlock_ioBundle_confOut[60:58]; // @[TileFull.scala 156:60]
  assign SBMux_C3_N23497_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C3_N23497_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C3_N23497_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C3_N23497_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C11_N23499_O_0_C_3_io_in = {SBMux_C11_N23499_O_0_C_3_io_in_hi,IN_CHANY_N32523_27}; // @[TileFull.scala 207:13]
  assign SBMux_C11_N23499_O_0_C_3_io_config = configBlock_ioBundle_confOut[63:61]; // @[TileFull.scala 156:60]
  assign SBMux_C11_N23499_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C11_N23499_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C11_N23499_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C11_N23499_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C19_N23501_O_0_C_3_io_in = {SBMux_C19_N23501_O_0_C_3_io_in_hi,IN_CHANY_N32515_19}; // @[TileFull.scala 207:13]
  assign SBMux_C19_N23501_O_0_C_3_io_config = configBlock_ioBundle_confOut[66:64]; // @[TileFull.scala 156:60]
  assign SBMux_C19_N23501_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C19_N23501_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C19_N23501_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C19_N23501_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C27_N23503_O_0_C_4_io_in = {SBMux_C27_N23503_O_0_C_4_io_in_hi,SBMux_C27_N23503_O_0_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C27_N23503_O_0_C_4_io_config = configBlock_ioBundle_confOut[69:67]; // @[TileFull.scala 156:60]
  assign SBMux_C27_N23503_O_0_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C27_N23503_O_0_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C27_N23503_O_0_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C27_N23503_O_0_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C35_N23505_O_0_C_3_io_in = {SBMux_C35_N23505_O_0_C_3_io_in_hi,IN_CHANY_N32507_11}; // @[TileFull.scala 207:13]
  assign SBMux_C35_N23505_O_0_C_3_io_config = configBlock_ioBundle_confOut[72:70]; // @[TileFull.scala 156:60]
  assign SBMux_C35_N23505_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C35_N23505_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C35_N23505_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C35_N23505_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C43_N23507_O_0_C_4_io_in = {SBMux_C43_N23507_O_0_C_4_io_in_hi,SBMux_C43_N23507_O_0_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C43_N23507_O_0_C_4_io_config = configBlock_ioBundle_confOut[75:73]; // @[TileFull.scala 156:60]
  assign SBMux_C43_N23507_O_0_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C43_N23507_O_0_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C43_N23507_O_0_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C43_N23507_O_0_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C51_N23509_O_0_C_2_io_in = {IN_CHANY_N32563_67,IN_CHANY_N32553_57}; // @[TileFull.scala 207:13]
  assign SBMux_C51_N23509_O_0_C_2_io_config = configBlock_ioBundle_confOut[77:76]; // @[TileFull.scala 156:60]
  assign SBMux_C51_N23509_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C51_N23509_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C51_N23509_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C51_N23509_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C59_N23511_O_0_C_3_io_in = {SBMux_C59_N23511_O_0_C_3_io_in_hi,IN_CHANY_N32497_1}; // @[TileFull.scala 207:13]
  assign SBMux_C59_N23511_O_0_C_3_io_config = configBlock_ioBundle_confOut[80:78]; // @[TileFull.scala 156:60]
  assign SBMux_C59_N23511_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C59_N23511_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C59_N23511_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C59_N23511_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C67_N23513_O_0_C_2_io_in = {IN_CHANY_N32593_97,IN_CHANY_N32575_79}; // @[TileFull.scala 207:13]
  assign SBMux_C67_N23513_O_0_C_2_io_config = configBlock_ioBundle_confOut[82:81]; // @[TileFull.scala 156:60]
  assign SBMux_C67_N23513_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C67_N23513_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C67_N23513_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C67_N23513_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C75_N23515_O_0_C_2_io_in = {IN_CHANY_N32591_95,IN_CHANY_N32571_75}; // @[TileFull.scala 207:13]
  assign SBMux_C75_N23515_O_0_C_2_io_config = configBlock_ioBundle_confOut[84:83]; // @[TileFull.scala 156:60]
  assign SBMux_C75_N23515_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C75_N23515_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C75_N23515_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C75_N23515_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C83_N23517_O_0_C_2_io_in = {IN_CHANY_N32603_107,IN_CHANY_N32539_43}; // @[TileFull.scala 207:13]
  assign SBMux_C83_N23517_O_0_C_2_io_config = configBlock_ioBundle_confOut[86:85]; // @[TileFull.scala 156:60]
  assign SBMux_C83_N23517_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C83_N23517_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C83_N23517_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C83_N23517_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C87_N23519_O_0_C_2_io_in = {IN_CHANY_N32581_85,IN_CHANY_N32511_15}; // @[TileFull.scala 207:13]
  assign SBMux_C87_N23519_O_0_C_2_io_config = configBlock_ioBundle_confOut[88:87]; // @[TileFull.scala 156:60]
  assign SBMux_C87_N23519_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C87_N23519_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C87_N23519_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C87_N23519_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C91_N23521_O_0_C_2_io_in = {IN_CHANY_N32585_89,IN_CHANY_N32497_1}; // @[TileFull.scala 207:13]
  assign SBMux_C91_N23521_O_0_C_2_io_config = configBlock_ioBundle_confOut[90:89]; // @[TileFull.scala 156:60]
  assign SBMux_C91_N23521_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C91_N23521_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C91_N23521_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C91_N23521_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C95_N23523_O_0_C_2_io_in = {IN_CHANY_N32601_105,IN_CHANY_N32519_23}; // @[TileFull.scala 207:13]
  assign SBMux_C95_N23523_O_0_C_2_io_config = configBlock_ioBundle_confOut[92:91]; // @[TileFull.scala 156:60]
  assign SBMux_C95_N23523_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C95_N23523_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C95_N23523_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C95_N23523_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C99_N23525_O_0_C_2_io_in = {IN_CHANY_N32579_83,IN_CHANY_N32547_51}; // @[TileFull.scala 207:13]
  assign SBMux_C99_N23525_O_0_C_2_io_config = configBlock_ioBundle_confOut[94:93]; // @[TileFull.scala 156:60]
  assign SBMux_C99_N23525_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C99_N23525_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C99_N23525_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C99_N23525_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C103_N23527_O_0_C_2_io_in = {IN_CHANY_N32583_87,IN_CHANY_N32525_29}; // @[TileFull.scala 207:13]
  assign SBMux_C103_N23527_O_0_C_2_io_config = configBlock_ioBundle_confOut[96:95]; // @[TileFull.scala 156:60]
  assign SBMux_C103_N23527_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C103_N23527_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C103_N23527_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C103_N23527_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C107_N23529_O_0_C_2_io_in = {IN_CHANY_N32597_101,IN_CHANY_N32517_21}; // @[TileFull.scala 207:13]
  assign SBMux_C107_N23529_O_0_C_2_io_config = configBlock_ioBundle_confOut[98:97]; // @[TileFull.scala 156:60]
  assign SBMux_C107_N23529_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C107_N23529_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C107_N23529_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C107_N23529_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C5_N23531_O_0_C_2_io_in = {IN_CHANY_N32567_71,IN_CHANY_N32549_53}; // @[TileFull.scala 207:13]
  assign SBMux_C5_N23531_O_0_C_2_io_config = configBlock_ioBundle_confOut[100:99]; // @[TileFull.scala 156:60]
  assign SBMux_C5_N23531_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C5_N23531_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C5_N23531_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C5_N23531_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C13_N23533_O_0_C_2_io_in = {IN_CHANY_N32577_81,IN_CHANY_N32503_7}; // @[TileFull.scala 207:13]
  assign SBMux_C13_N23533_O_0_C_2_io_config = configBlock_ioBundle_confOut[102:101]; // @[TileFull.scala 156:60]
  assign SBMux_C13_N23533_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C13_N23533_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C13_N23533_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C13_N23533_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C21_N23535_O_0_C_3_io_in = {SBMux_C21_N23535_O_0_C_3_io_in_hi,IN_CHANY_N32547_51}; // @[TileFull.scala 207:13]
  assign SBMux_C21_N23535_O_0_C_3_io_config = configBlock_ioBundle_confOut[105:103]; // @[TileFull.scala 156:60]
  assign SBMux_C21_N23535_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C21_N23535_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C21_N23535_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C21_N23535_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C29_N23537_O_0_C_2_io_in = {IN_CHANY_N32579_83,IN_CHANY_N32557_61}; // @[TileFull.scala 207:13]
  assign SBMux_C29_N23537_O_0_C_2_io_config = configBlock_ioBundle_confOut[107:106]; // @[TileFull.scala 156:60]
  assign SBMux_C29_N23537_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C29_N23537_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C29_N23537_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C29_N23537_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C37_N23539_O_0_C_3_io_in = {SBMux_C37_N23539_O_0_C_3_io_in_hi,IN_CHANY_N32527_31}; // @[TileFull.scala 207:13]
  assign SBMux_C37_N23539_O_0_C_3_io_config = configBlock_ioBundle_confOut[110:108]; // @[TileFull.scala 156:60]
  assign SBMux_C37_N23539_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C37_N23539_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C37_N23539_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C37_N23539_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C45_N23541_O_0_C_2_io_in = {IN_CHANY_N32569_73,IN_CHANY_N32545_49}; // @[TileFull.scala 207:13]
  assign SBMux_C45_N23541_O_0_C_2_io_config = configBlock_ioBundle_confOut[112:111]; // @[TileFull.scala 156:60]
  assign SBMux_C45_N23541_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C45_N23541_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C45_N23541_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C45_N23541_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C53_N23543_O_0_C_3_io_in = {SBMux_C25_N23469_O_0_C_3_io_in_hi,IN_CHANY_N32521_25}; // @[TileFull.scala 207:13]
  assign SBMux_C53_N23543_O_0_C_3_io_config = configBlock_ioBundle_confOut[115:113]; // @[TileFull.scala 156:60]
  assign SBMux_C53_N23543_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C53_N23543_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C53_N23543_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C53_N23543_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C61_N23545_O_0_C_3_io_in = {SBMux_C61_N23545_O_0_C_3_io_in_hi,IN_CHANY_N32519_23}; // @[TileFull.scala 207:13]
  assign SBMux_C61_N23545_O_0_C_3_io_config = configBlock_ioBundle_confOut[118:116]; // @[TileFull.scala 156:60]
  assign SBMux_C61_N23545_O_0_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C61_N23545_O_0_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C61_N23545_O_0_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C61_N23545_O_0_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C69_N23547_O_0_C_2_io_in = {IN_CHANY_N32579_83,IN_CHANY_N32569_73}; // @[TileFull.scala 207:13]
  assign SBMux_C69_N23547_O_0_C_2_io_config = configBlock_ioBundle_confOut[120:119]; // @[TileFull.scala 156:60]
  assign SBMux_C69_N23547_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C69_N23547_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C69_N23547_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C69_N23547_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C77_N23549_O_0_C_2_io_in = {IN_CHANY_N32587_91,IN_CHANY_N32573_77}; // @[TileFull.scala 207:13]
  assign SBMux_C77_N23549_O_0_C_2_io_config = configBlock_ioBundle_confOut[122:121]; // @[TileFull.scala 156:60]
  assign SBMux_C77_N23549_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C77_N23549_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C77_N23549_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C77_N23549_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C85_N23551_O_0_C_2_io_in = {IN_CHANY_N32589_93,IN_CHANY_N32557_61}; // @[TileFull.scala 207:13]
  assign SBMux_C85_N23551_O_0_C_2_io_config = configBlock_ioBundle_confOut[124:123]; // @[TileFull.scala 156:60]
  assign SBMux_C85_N23551_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C85_N23551_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C85_N23551_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C85_N23551_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C89_N23553_O_0_C_2_io_in = {IN_CHANY_N32595_99,IN_CHANY_N32537_41}; // @[TileFull.scala 207:13]
  assign SBMux_C89_N23553_O_0_C_2_io_config = configBlock_ioBundle_confOut[126:125]; // @[TileFull.scala 156:60]
  assign SBMux_C89_N23553_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C89_N23553_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C89_N23553_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C89_N23553_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C93_N23555_O_0_C_2_io_in = {IN_CHANY_N32593_97,IN_CHANY_N32551_55}; // @[TileFull.scala 207:13]
  assign SBMux_C93_N23555_O_0_C_2_io_config = configBlock_ioBundle_confOut[128:127]; // @[TileFull.scala 156:60]
  assign SBMux_C93_N23555_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C93_N23555_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C93_N23555_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C93_N23555_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C97_N23557_O_0_C_2_io_in = {IN_CHANY_N32587_91,IN_CHANY_N32543_47}; // @[TileFull.scala 207:13]
  assign SBMux_C97_N23557_O_0_C_2_io_config = configBlock_ioBundle_confOut[130:129]; // @[TileFull.scala 156:60]
  assign SBMux_C97_N23557_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C97_N23557_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C97_N23557_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C97_N23557_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C101_N23559_O_0_C_2_io_in = {IN_CHANY_N32599_103,IN_CHANY_N32545_49}; // @[TileFull.scala 207:13]
  assign SBMux_C101_N23559_O_0_C_2_io_config = configBlock_ioBundle_confOut[132:131]; // @[TileFull.scala 156:60]
  assign SBMux_C101_N23559_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C101_N23559_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C101_N23559_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C101_N23559_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C105_N23561_O_0_C_2_io_in = {IN_CHANY_N32591_95,IN_CHANY_N32561_65}; // @[TileFull.scala 207:13]
  assign SBMux_C105_N23561_O_0_C_2_io_config = configBlock_ioBundle_confOut[134:133]; // @[TileFull.scala 156:60]
  assign SBMux_C105_N23561_O_0_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C105_N23561_O_0_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C105_N23561_O_0_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C105_N23561_O_0_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C0_N32496_O_2_C_3_io_in = {SBMux_C0_N32496_O_2_C_3_io_in_hi,SBMux_C0_N32496_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C0_N32496_O_2_C_3_io_config = configBlock_ioBundle_confOut[137:135]; // @[TileFull.scala 156:60]
  assign SBMux_C0_N32496_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C0_N32496_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C0_N32496_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C0_N32496_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C2_N32498_O_2_C_3_io_in = {SBMux_C2_N32498_O_2_C_3_io_in_hi,SBMux_C2_N32498_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C2_N32498_O_2_C_3_io_config = configBlock_ioBundle_confOut[140:138]; // @[TileFull.scala 156:60]
  assign SBMux_C2_N32498_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C2_N32498_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C2_N32498_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C2_N32498_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C4_N32500_O_2_C_3_io_in = {SBMux_C4_N32500_O_2_C_3_io_in_hi,SBMux_C4_N32500_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C4_N32500_O_2_C_3_io_config = configBlock_ioBundle_confOut[143:141]; // @[TileFull.scala 156:60]
  assign SBMux_C4_N32500_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C4_N32500_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C4_N32500_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C4_N32500_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C6_N32502_O_2_C_4_io_in = {SBMux_C6_N32502_O_2_C_4_io_in_hi,SBMux_C6_N32502_O_2_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C6_N32502_O_2_C_4_io_config = configBlock_ioBundle_confOut[146:144]; // @[TileFull.scala 156:60]
  assign SBMux_C6_N32502_O_2_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C6_N32502_O_2_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C6_N32502_O_2_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C6_N32502_O_2_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C8_N32504_O_2_C_3_io_in = {SBMux_C8_N32504_O_2_C_3_io_in_hi,SBMux_C8_N32504_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C8_N32504_O_2_C_3_io_config = configBlock_ioBundle_confOut[149:147]; // @[TileFull.scala 156:60]
  assign SBMux_C8_N32504_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C8_N32504_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C8_N32504_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C8_N32504_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C10_N32506_O_2_C_4_io_in = {SBMux_C10_N32506_O_2_C_4_io_in_hi,SBMux_C10_N32506_O_2_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C10_N32506_O_2_C_4_io_config = configBlock_ioBundle_confOut[152:150]; // @[TileFull.scala 156:60]
  assign SBMux_C10_N32506_O_2_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C10_N32506_O_2_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C10_N32506_O_2_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C10_N32506_O_2_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C12_N32508_O_2_C_3_io_in = {SBMux_C12_N32508_O_2_C_3_io_in_hi,SBMux_C12_N32508_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C12_N32508_O_2_C_3_io_config = configBlock_ioBundle_confOut[155:153]; // @[TileFull.scala 156:60]
  assign SBMux_C12_N32508_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C12_N32508_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C12_N32508_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C12_N32508_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C14_N32510_O_2_C_4_io_in = {SBMux_C14_N32510_O_2_C_4_io_in_hi,SBMux_C14_N32510_O_2_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C14_N32510_O_2_C_4_io_config = configBlock_ioBundle_confOut[158:156]; // @[TileFull.scala 156:60]
  assign SBMux_C14_N32510_O_2_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C14_N32510_O_2_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C14_N32510_O_2_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C14_N32510_O_2_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C16_N32512_O_2_C_3_io_in = {SBMux_C16_N32512_O_2_C_3_io_in_hi,SBMux_C16_N32512_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C16_N32512_O_2_C_3_io_config = configBlock_ioBundle_confOut[161:159]; // @[TileFull.scala 156:60]
  assign SBMux_C16_N32512_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C16_N32512_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C16_N32512_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C16_N32512_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C18_N32514_O_2_C_4_io_in = {SBMux_C18_N32514_O_2_C_4_io_in_hi,SBMux_C18_N32514_O_2_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C18_N32514_O_2_C_4_io_config = configBlock_ioBundle_confOut[164:162]; // @[TileFull.scala 156:60]
  assign SBMux_C18_N32514_O_2_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C18_N32514_O_2_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C18_N32514_O_2_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C18_N32514_O_2_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C20_N32516_O_2_C_4_io_in = {SBMux_C20_N32516_O_2_C_4_io_in_hi,SBMux_C20_N32516_O_2_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C20_N32516_O_2_C_4_io_config = configBlock_ioBundle_confOut[167:165]; // @[TileFull.scala 156:60]
  assign SBMux_C20_N32516_O_2_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C20_N32516_O_2_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C20_N32516_O_2_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C20_N32516_O_2_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C22_N32518_O_2_C_3_io_in = {SBMux_C22_N32518_O_2_C_3_io_in_hi,SBMux_C22_N32518_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C22_N32518_O_2_C_3_io_config = configBlock_ioBundle_confOut[170:168]; // @[TileFull.scala 156:60]
  assign SBMux_C22_N32518_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C22_N32518_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C22_N32518_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C22_N32518_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C24_N32520_O_2_C_2_io_in = {SBMux_C24_N32520_O_2_C_2_io_in_hi,SBMux_C24_N32520_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C24_N32520_O_2_C_2_io_config = configBlock_ioBundle_confOut[172:171]; // @[TileFull.scala 156:60]
  assign SBMux_C24_N32520_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C24_N32520_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C24_N32520_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C24_N32520_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C26_N32522_O_2_C_3_io_in = {SBMux_C26_N32522_O_2_C_3_io_in_hi,SBMux_C26_N32522_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C26_N32522_O_2_C_3_io_config = configBlock_ioBundle_confOut[175:173]; // @[TileFull.scala 156:60]
  assign SBMux_C26_N32522_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C26_N32522_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C26_N32522_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C26_N32522_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C28_N32524_O_2_C_2_io_in = {SBMux_C28_N32524_O_2_C_2_io_in_hi,SBMux_C28_N32524_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C28_N32524_O_2_C_2_io_config = configBlock_ioBundle_confOut[177:176]; // @[TileFull.scala 156:60]
  assign SBMux_C28_N32524_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C28_N32524_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C28_N32524_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C28_N32524_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C30_N32526_O_2_C_2_io_in = {SBMux_C30_N32526_O_2_C_2_io_in_hi,SBMux_C30_N32526_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C30_N32526_O_2_C_2_io_config = configBlock_ioBundle_confOut[179:178]; // @[TileFull.scala 156:60]
  assign SBMux_C30_N32526_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C30_N32526_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C30_N32526_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C30_N32526_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C32_N32528_O_2_C_4_io_in = {SBMux_C32_N32528_O_2_C_4_io_in_hi,SBMux_C32_N32528_O_2_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C32_N32528_O_2_C_4_io_config = configBlock_ioBundle_confOut[182:180]; // @[TileFull.scala 156:60]
  assign SBMux_C32_N32528_O_2_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C32_N32528_O_2_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C32_N32528_O_2_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C32_N32528_O_2_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C34_N32530_O_2_C_3_io_in = {SBMux_C34_N32530_O_2_C_3_io_in_hi,SBMux_C34_N32530_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C34_N32530_O_2_C_3_io_config = configBlock_ioBundle_confOut[185:183]; // @[TileFull.scala 156:60]
  assign SBMux_C34_N32530_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C34_N32530_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C34_N32530_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C34_N32530_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C36_N32532_O_2_C_3_io_in = {SBMux_C36_N32532_O_2_C_3_io_in_hi,SBMux_C36_N32532_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C36_N32532_O_2_C_3_io_config = configBlock_ioBundle_confOut[188:186]; // @[TileFull.scala 156:60]
  assign SBMux_C36_N32532_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C36_N32532_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C36_N32532_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C36_N32532_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C38_N32534_O_2_C_4_io_in = {SBMux_C38_N32534_O_2_C_4_io_in_hi,SBMux_C38_N32534_O_2_C_4_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C38_N32534_O_2_C_4_io_config = configBlock_ioBundle_confOut[191:189]; // @[TileFull.scala 156:60]
  assign SBMux_C38_N32534_O_2_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C38_N32534_O_2_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C38_N32534_O_2_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C38_N32534_O_2_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C40_N32536_O_2_C_2_io_in = {SBMux_C40_N32536_O_2_C_2_io_in_hi,SBMux_C40_N32536_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C40_N32536_O_2_C_2_io_config = configBlock_ioBundle_confOut[193:192]; // @[TileFull.scala 156:60]
  assign SBMux_C40_N32536_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C40_N32536_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C40_N32536_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C40_N32536_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C42_N32538_O_2_C_3_io_in = {SBMux_C42_N32538_O_2_C_3_io_in_hi,SBMux_C42_N32538_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C42_N32538_O_2_C_3_io_config = configBlock_ioBundle_confOut[196:194]; // @[TileFull.scala 156:60]
  assign SBMux_C42_N32538_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C42_N32538_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C42_N32538_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C42_N32538_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C44_N32540_O_2_C_3_io_in = {SBMux_C44_N32540_O_2_C_3_io_in_hi,SBMux_C44_N32540_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C44_N32540_O_2_C_3_io_config = configBlock_ioBundle_confOut[199:197]; // @[TileFull.scala 156:60]
  assign SBMux_C44_N32540_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C44_N32540_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C44_N32540_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C44_N32540_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C46_N32542_O_2_C_3_io_in = {SBMux_C46_N32542_O_2_C_3_io_in_hi,SBMux_C46_N32542_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C46_N32542_O_2_C_3_io_config = configBlock_ioBundle_confOut[202:200]; // @[TileFull.scala 156:60]
  assign SBMux_C46_N32542_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C46_N32542_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C46_N32542_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C46_N32542_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C48_N32544_O_2_C_3_io_in = {SBMux_C48_N32544_O_2_C_3_io_in_hi,SBMux_C48_N32544_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C48_N32544_O_2_C_3_io_config = configBlock_ioBundle_confOut[205:203]; // @[TileFull.scala 156:60]
  assign SBMux_C48_N32544_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C48_N32544_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C48_N32544_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C48_N32544_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C50_N32546_O_2_C_3_io_in = {SBMux_C50_N32546_O_2_C_3_io_in_hi,SBMux_C50_N32546_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C50_N32546_O_2_C_3_io_config = configBlock_ioBundle_confOut[208:206]; // @[TileFull.scala 156:60]
  assign SBMux_C50_N32546_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C50_N32546_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C50_N32546_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C50_N32546_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C52_N32548_O_2_C_3_io_in = {SBMux_C52_N32548_O_2_C_3_io_in_hi,SBMux_C52_N32548_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C52_N32548_O_2_C_3_io_config = configBlock_ioBundle_confOut[211:209]; // @[TileFull.scala 156:60]
  assign SBMux_C52_N32548_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C52_N32548_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C52_N32548_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C52_N32548_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C54_N32550_O_2_C_2_io_in = {SBMux_C54_N32550_O_2_C_2_io_in_hi,SBMux_C54_N32550_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C54_N32550_O_2_C_2_io_config = configBlock_ioBundle_confOut[213:212]; // @[TileFull.scala 156:60]
  assign SBMux_C54_N32550_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C54_N32550_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C54_N32550_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C54_N32550_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C56_N32552_O_2_C_3_io_in = {SBMux_C56_N32552_O_2_C_3_io_in_hi,SBMux_C56_N32552_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C56_N32552_O_2_C_3_io_config = configBlock_ioBundle_confOut[216:214]; // @[TileFull.scala 156:60]
  assign SBMux_C56_N32552_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C56_N32552_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C56_N32552_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C56_N32552_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C58_N32554_O_2_C_2_io_in = {SBMux_C58_N32554_O_2_C_2_io_in_hi,SBMux_C58_N32554_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C58_N32554_O_2_C_2_io_config = configBlock_ioBundle_confOut[218:217]; // @[TileFull.scala 156:60]
  assign SBMux_C58_N32554_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C58_N32554_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C58_N32554_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C58_N32554_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C60_N32556_O_2_C_3_io_in = {SBMux_C60_N32556_O_2_C_3_io_in_hi,SBMux_C60_N32556_O_2_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C60_N32556_O_2_C_3_io_config = configBlock_ioBundle_confOut[221:219]; // @[TileFull.scala 156:60]
  assign SBMux_C60_N32556_O_2_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C60_N32556_O_2_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C60_N32556_O_2_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C60_N32556_O_2_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C62_N32558_O_1_C_3_io_in = {SBMux_C62_N32558_O_1_C_3_io_in_hi,SBMux_C62_N32558_O_1_C_3_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C62_N32558_O_1_C_3_io_config = configBlock_ioBundle_confOut[224:222]; // @[TileFull.scala 156:60]
  assign SBMux_C62_N32558_O_1_C_3_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C62_N32558_O_1_C_3_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C62_N32558_O_1_C_3_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C62_N32558_O_1_C_3_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C64_N32560_O_1_C_2_io_in = {SBMux_C64_N32560_O_1_C_2_io_in_hi,IN_OPIN_N21952_48}; // @[TileFull.scala 207:13]
  assign SBMux_C64_N32560_O_1_C_2_io_config = configBlock_ioBundle_confOut[226:225]; // @[TileFull.scala 156:60]
  assign SBMux_C64_N32560_O_1_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C64_N32560_O_1_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C64_N32560_O_1_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C64_N32560_O_1_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C66_N32562_O_4_C_2_io_in = {SBMux_C66_N32562_O_4_C_2_io_in_hi,SBMux_C66_N32562_O_4_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C66_N32562_O_4_C_2_io_config = configBlock_ioBundle_confOut[229:227]; // @[TileFull.scala 156:60]
  assign SBMux_C66_N32562_O_4_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C66_N32562_O_4_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C66_N32562_O_4_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C66_N32562_O_4_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C68_N32564_O_4_C_2_io_in = {SBMux_C68_N32564_O_4_C_2_io_in_hi,SBMux_C68_N32564_O_4_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C68_N32564_O_4_C_2_io_config = configBlock_ioBundle_confOut[232:230]; // @[TileFull.scala 156:60]
  assign SBMux_C68_N32564_O_4_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C68_N32564_O_4_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C68_N32564_O_4_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C68_N32564_O_4_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C70_N32566_O_4_C_2_io_in = {SBMux_C70_N32566_O_4_C_2_io_in_hi,SBMux_C70_N32566_O_4_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C70_N32566_O_4_C_2_io_config = configBlock_ioBundle_confOut[235:233]; // @[TileFull.scala 156:60]
  assign SBMux_C70_N32566_O_4_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C70_N32566_O_4_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C70_N32566_O_4_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C70_N32566_O_4_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C72_N32568_O_4_C_2_io_in = {SBMux_C72_N32568_O_4_C_2_io_in_hi,SBMux_C72_N32568_O_4_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C72_N32568_O_4_C_2_io_config = configBlock_ioBundle_confOut[238:236]; // @[TileFull.scala 156:60]
  assign SBMux_C72_N32568_O_4_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C72_N32568_O_4_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C72_N32568_O_4_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C72_N32568_O_4_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C74_N32570_O_4_C_2_io_in = {SBMux_C74_N32570_O_4_C_2_io_in_hi,SBMux_C74_N32570_O_4_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C74_N32570_O_4_C_2_io_config = configBlock_ioBundle_confOut[241:239]; // @[TileFull.scala 156:60]
  assign SBMux_C74_N32570_O_4_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C74_N32570_O_4_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C74_N32570_O_4_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C74_N32570_O_4_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C76_N32572_O_4_C_2_io_in = {SBMux_C76_N32572_O_4_C_2_io_in_hi,SBMux_C76_N32572_O_4_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C76_N32572_O_4_C_2_io_config = configBlock_ioBundle_confOut[244:242]; // @[TileFull.scala 156:60]
  assign SBMux_C76_N32572_O_4_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C76_N32572_O_4_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C76_N32572_O_4_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C76_N32572_O_4_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C78_N32574_O_4_C_2_io_in = {SBMux_C78_N32574_O_4_C_2_io_in_hi,SBMux_C78_N32574_O_4_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C78_N32574_O_4_C_2_io_config = configBlock_ioBundle_confOut[247:245]; // @[TileFull.scala 156:60]
  assign SBMux_C78_N32574_O_4_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C78_N32574_O_4_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C78_N32574_O_4_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C78_N32574_O_4_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C80_N32576_O_4_C_2_io_in = {SBMux_C80_N32576_O_4_C_2_io_in_hi,SBMux_C80_N32576_O_4_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C80_N32576_O_4_C_2_io_config = configBlock_ioBundle_confOut[250:248]; // @[TileFull.scala 156:60]
  assign SBMux_C80_N32576_O_4_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C80_N32576_O_4_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C80_N32576_O_4_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C80_N32576_O_4_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C82_N32578_O_3_C_2_io_in = {SBMux_C82_N32578_O_3_C_2_io_in_hi,SBMux_C82_N32578_O_3_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C82_N32578_O_3_C_2_io_config = configBlock_ioBundle_confOut[253:251]; // @[TileFull.scala 156:60]
  assign SBMux_C82_N32578_O_3_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C82_N32578_O_3_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C82_N32578_O_3_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C82_N32578_O_3_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C84_N32580_O_3_C_2_io_in = {SBMux_C84_N32580_O_3_C_2_io_in_hi,SBMux_C84_N32580_O_3_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C84_N32580_O_3_C_2_io_config = configBlock_ioBundle_confOut[256:254]; // @[TileFull.scala 156:60]
  assign SBMux_C84_N32580_O_3_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C84_N32580_O_3_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C84_N32580_O_3_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C84_N32580_O_3_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C86_N32582_O_3_C_2_io_in = {SBMux_C86_N32582_O_3_C_2_io_in_hi,SBMux_C86_N32582_O_3_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C86_N32582_O_3_C_2_io_config = configBlock_ioBundle_confOut[259:257]; // @[TileFull.scala 156:60]
  assign SBMux_C86_N32582_O_3_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C86_N32582_O_3_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C86_N32582_O_3_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C86_N32582_O_3_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C88_N32584_O_3_C_2_io_in = {SBMux_C88_N32584_O_3_C_2_io_in_hi,SBMux_C88_N32584_O_3_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C88_N32584_O_3_C_2_io_config = configBlock_ioBundle_confOut[262:260]; // @[TileFull.scala 156:60]
  assign SBMux_C88_N32584_O_3_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C88_N32584_O_3_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C88_N32584_O_3_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C88_N32584_O_3_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C90_N32586_O_3_C_2_io_in = {SBMux_C90_N32586_O_3_C_2_io_in_hi,SBMux_C90_N32586_O_3_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C90_N32586_O_3_C_2_io_config = configBlock_ioBundle_confOut[265:263]; // @[TileFull.scala 156:60]
  assign SBMux_C90_N32586_O_3_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C90_N32586_O_3_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C90_N32586_O_3_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C90_N32586_O_3_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C92_N32588_O_3_C_2_io_in = {SBMux_C92_N32588_O_3_C_2_io_in_hi,SBMux_C92_N32588_O_3_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C92_N32588_O_3_C_2_io_config = configBlock_ioBundle_confOut[268:266]; // @[TileFull.scala 156:60]
  assign SBMux_C92_N32588_O_3_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C92_N32588_O_3_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C92_N32588_O_3_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C92_N32588_O_3_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C94_N32590_O_2_C_2_io_in = {SBMux_C94_N32590_O_2_C_2_io_in_hi,SBMux_C94_N32590_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C94_N32590_O_2_C_2_io_config = configBlock_ioBundle_confOut[270:269]; // @[TileFull.scala 156:60]
  assign SBMux_C94_N32590_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C94_N32590_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C94_N32590_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C94_N32590_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C96_N32592_O_2_C_2_io_in = {SBMux_C96_N32592_O_2_C_2_io_in_hi,SBMux_C96_N32592_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C96_N32592_O_2_C_2_io_config = configBlock_ioBundle_confOut[272:271]; // @[TileFull.scala 156:60]
  assign SBMux_C96_N32592_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C96_N32592_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C96_N32592_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C96_N32592_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C98_N32594_O_2_C_2_io_in = {SBMux_C98_N32594_O_2_C_2_io_in_hi,SBMux_C98_N32594_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C98_N32594_O_2_C_2_io_config = configBlock_ioBundle_confOut[274:273]; // @[TileFull.scala 156:60]
  assign SBMux_C98_N32594_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C98_N32594_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C98_N32594_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C98_N32594_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C100_N32596_O_2_C_2_io_in = {SBMux_C100_N32596_O_2_C_2_io_in_hi,SBMux_C100_N32596_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C100_N32596_O_2_C_2_io_config = configBlock_ioBundle_confOut[276:275]; // @[TileFull.scala 156:60]
  assign SBMux_C100_N32596_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C100_N32596_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C100_N32596_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C100_N32596_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C102_N32598_O_2_C_2_io_in = {SBMux_C102_N32598_O_2_C_2_io_in_hi,SBMux_C102_N32598_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C102_N32598_O_2_C_2_io_config = configBlock_ioBundle_confOut[278:277]; // @[TileFull.scala 156:60]
  assign SBMux_C102_N32598_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C102_N32598_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C102_N32598_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C102_N32598_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C104_N32600_O_2_C_2_io_in = {SBMux_C104_N32600_O_2_C_2_io_in_hi,SBMux_C104_N32600_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C104_N32600_O_2_C_2_io_config = configBlock_ioBundle_confOut[280:279]; // @[TileFull.scala 156:60]
  assign SBMux_C104_N32600_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C104_N32600_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C104_N32600_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C104_N32600_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
  assign SBMux_C106_N32602_O_2_C_2_io_in = {SBMux_C36_N32532_O_2_C_3_io_in_hi_hi,SBMux_C106_N32602_O_2_C_2_io_in_lo}; // @[TileFull.scala 207:13]
  assign SBMux_C106_N32602_O_2_C_2_io_config = configBlock_ioBundle_confOut[282:281]; // @[TileFull.scala 156:60]
  assign SBMux_C106_N32602_O_2_C_2_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 160:28]
  assign SBMux_C106_N32602_O_2_C_2_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 163:27]
  assign SBMux_C106_N32602_O_2_C_2_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 161:26]
  assign SBMux_C106_N32602_O_2_C_2_io_arst = ctrlSignals_arst; // @[TileFull.scala 162:23]
endmodule
