/afs/ece.cmu.edu/project/km_group/.vol9/asap7/asap7sc7p5t_28/techlef_misc/asap7_tech_4x_201209_mod.lef