module AluMul(
  input         clock,
  input         reset,
  input  [15:0] io_i0,
  input  [15:0] io_i1,
  input  [31:0] io_ib32,
  input  [7:0]  io_ctrl,
  output [15:0] io_q,
  input  [31:0] io_config,
  input         io_gndOuts,
  input         io_clkEnb,
  input         io_loopBreak
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  _i0FF_T = ~io_clkEnb; // @[CLBlut4N10Mul.scala 100:44]
  reg [15:0] i0FF; // @[Reg.scala 28:20]
  reg [15:0] i1FF; // @[Reg.scala 28:20]
  reg [31:0] ib32FF; // @[Reg.scala 28:20]
  wire [15:0] in0 = io_config[0] ? io_i0 : i0FF; // @[CLBlut4N10Mul.scala 104:44]
  wire [15:0] in1 = io_config[1] ? io_i1 : i1FF; // @[CLBlut4N10Mul.scala 105:44]
  wire [31:0] ib32 = io_config[2] ? io_ib32 : ib32FF; // @[CLBlut4N10Mul.scala 106:49]
  wire [15:0] _add_T_2 = $signed(in0) + $signed(in1); // @[CLBlut4N10Mul.scala 108:17]
  wire [31:0] _GEN_4 = {{16{_add_T_2[15]}},_add_T_2}; // @[CLBlut4N10Mul.scala 108:23]
  wire [31:0] add = $signed(_GEN_4) + $signed(ib32); // @[CLBlut4N10Mul.scala 108:23]
  wire [31:0] mul16 = $signed(in0) * $signed(in1); // @[CLBlut4N10Mul.scala 110:16]
  wire [15:0] mux_lo = io_ctrl[3] ? $signed(in1) : $signed(in0); // @[Cat.scala 31:58]
  wire [31:0] mux = {16'h0,mux_lo}; // @[CLBlut4N10Mul.scala 111:60]
  wire [1:0] _accVal_T_2 = {io_config[4],io_config[3]}; // @[Cat.scala 31:58]
  reg [31:0] accFF_r; // @[Reg.scala 28:20]
  wire [31:0] accVal = _accVal_T_2 == 2'h2 ? $signed(accFF_r) : $signed(32'sh0); // @[CLBlut4N10Mul.scala 113:19]
  wire [31:0] _mac_T_2 = $signed(mul16) + $signed(ib32); // @[CLBlut4N10Mul.scala 114:19]
  wire [31:0] mac = $signed(_mac_T_2) + $signed(accVal); // @[CLBlut4N10Mul.scala 114:26]
  wire [31:0] _combOut_T_4 = 2'h1 == _accVal_T_2 ? $signed(mul16) : $signed(add); // @[Mux.scala 81:58]
  wire [31:0] _combOut_T_6 = 2'h2 == _accVal_T_2 ? $signed(mac) : $signed(_combOut_T_4); // @[Mux.scala 81:58]
  wire [31:0] combOut = 2'h3 == _accVal_T_2 ? $signed(mux) : $signed(_combOut_T_6); // @[Mux.scala 81:58]
  wire  _accFF_T_4 = io_ctrl[1] & _i0FF_T; // @[CLBlut4N10Mul.scala 117:69]
  wire [31:0] _out_T_3 = io_config[7] | io_loopBreak ? $signed(accFF_r) : $signed(combOut); // @[CLBlut4N10Mul.scala 120:83]
  wire [31:0] out = io_gndOuts ? 32'h0 : _out_T_3; // @[CLBlut4N10Mul.scala 120:16]
  assign io_q = io_ctrl[2] ? out[31:16] : out[15:0]; // @[CLBlut4N10Mul.scala 122:14]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      i0FF <= 16'h0; // @[Reg.scala 28:20]
    end else if (_i0FF_T) begin // @[Reg.scala 29:18]
      i0FF <= io_i0; // @[Reg.scala 29:22]
    end
    if (reset) begin // @[Reg.scala 28:20]
      i1FF <= 16'h0; // @[Reg.scala 28:20]
    end else if (_i0FF_T) begin // @[Reg.scala 29:18]
      i1FF <= io_i1; // @[Reg.scala 29:22]
    end
    if (reset) begin // @[Reg.scala 28:20]
      ib32FF <= 32'h0; // @[Reg.scala 28:20]
    end else if (_i0FF_T) begin // @[Reg.scala 29:18]
      ib32FF <= io_ib32; // @[Reg.scala 29:22]
    end
    if (reset) begin // @[Reg.scala 28:20]
      accFF_r <= 32'sh0; // @[Reg.scala 28:20]
    end else if (_accFF_T_4) begin // @[Reg.scala 29:18]
      if (io_ctrl[0]) begin // @[CLBlut4N10Mul.scala 117:25]
        accFF_r <= 32'sh0;
      end else if (2'h3 == _accVal_T_2) begin // @[Mux.scala 81:58]
        accFF_r <= mux;
      end else begin
        accFF_r <= _combOut_T_6;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i0FF = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  i1FF = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  ib32FF = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  accFF_r = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Ble4(
  input         clock,
  input         reset,
  input  [19:0] io_config,
  input         io_in_0,
  input         io_in_1,
  input         io_in_2,
  input         io_in_3,
  output        io_outR,
  output        io_outT,
  input         io_gndOuts,
  input         io_clkEnb,
  input         io_loopBreak
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] lut_in; // @[CLBlut4N10Clb.scala 76:27]
  wire [3:0] lut_sel; // @[CLBlut4N10Clb.scala 76:27]
  wire  lut_o; // @[CLBlut4N10Clb.scala 76:27]
  wire [1:0] lut_io_sel_lo = {io_in_1,io_in_0}; // @[CLBlut4N10Clb.scala 78:23]
  wire [1:0] lut_io_sel_hi = {io_in_3,io_in_2}; // @[CLBlut4N10Clb.scala 78:23]
  wire  _bleFF_T = ~io_clkEnb; // @[CLBlut4N10Clb.scala 80:48]
  reg  bleFF; // @[Reg.scala 28:20]
  wire  _io_outR_T_1 = ~io_loopBreak; // @[CLBlut4N10Clb.scala 83:34]
  wire  _io_outR_T_3 = io_config[16] & ~io_loopBreak ? lut_o : bleFF; // @[CLBlut4N10Clb.scala 83:17]
  wire  _io_outR_T_4 = ~io_gndOuts; // @[CLBlut4N10Clb.scala 83:68]
  wire  _io_outT_T_3 = io_config[17] & _io_outR_T_1 ? lut_o : bleFF; // @[CLBlut4N10Clb.scala 84:17]
  Mux16C lut ( // @[CLBlut4N10Clb.scala 76:27]
    .in(lut_in),
    .sel(lut_sel),
    .o(lut_o)
  );
  assign io_outR = _io_outR_T_3 & ~io_gndOuts; // @[CLBlut4N10Clb.scala 83:66]
  assign io_outT = _io_outT_T_3 & _io_outR_T_4; // @[CLBlut4N10Clb.scala 84:66]
  assign lut_in = io_config[15:0]; // @[CLBlut4N10Clb.scala 77:25]
  assign lut_sel = {lut_io_sel_hi,lut_io_sel_lo}; // @[CLBlut4N10Clb.scala 78:23]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      bleFF <= 1'h0; // @[Reg.scala 28:20]
    end else if (_bleFF_T) begin // @[Reg.scala 29:18]
      bleFF <= lut_o; // @[Reg.scala 29:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bleFF = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLBlut4N10Mul(
  input          IPIN_0,
  input          IPIN_1,
  input          IPIN_2,
  input          IPIN_3,
  input          IPIN_4,
  input          IPIN_5,
  input          IPIN_6,
  input          IPIN_7,
  input          IPIN_8,
  input          IPIN_9,
  input          IPIN_10,
  input          IPIN_11,
  input          IPIN_12,
  input          IPIN_13,
  input          IPIN_14,
  input          IPIN_15,
  input          IPIN_16,
  input          IPIN_17,
  input          IPIN_18,
  input          IPIN_19,
  input          IPIN_20,
  input          IPIN_21,
  input          IPIN_22,
  input          IPIN_23,
  input          IPIN_24,
  input          IPIN_25,
  input          IPIN_26,
  input          IPIN_27,
  input          IPIN_28,
  input          IPIN_29,
  input          IPIN_30,
  input          IPIN_31,
  input          IPIN_32,
  input          IPIN_33,
  input          IPIN_34,
  input          IPIN_35,
  input          IPIN_36,
  input          IPIN_37,
  input          IPIN_38,
  input          IPIN_39,
  input          IPIN_40,
  input          IPIN_41,
  input          IPIN_42,
  input          IPIN_43,
  input          IPIN_44,
  input          IPIN_45,
  input          IPIN_46,
  input          IPIN_47,
  input          IPIN_48,
  input          IPIN_49,
  input          IPIN_50,
  input          IPIN_51,
  input          IPIN_52,
  input          IPIN_53,
  input          IPIN_54,
  input          IPIN_55,
  input          IPIN_56,
  input          IPIN_57,
  input          IPIN_58,
  input          IPIN_59,
  input          IPIN_60,
  input          IPIN_61,
  input          IPIN_62,
  input          IPIN_63,
  input          IPIN_64,
  input          IPIN_65,
  input          IPIN_66,
  input          IPIN_67,
  input          IPIN_68,
  input          IPIN_69,
  input          IPIN_70,
  input          IPIN_71,
  output         OPIN_73,
  output         OPIN_74,
  output         OPIN_75,
  output         OPIN_76,
  output         OPIN_77,
  output         OPIN_78,
  output         OPIN_79,
  output         OPIN_80,
  output         OPIN_81,
  output         OPIN_82,
  output         OPIN_83,
  output         OPIN_84,
  output         OPIN_85,
  output         OPIN_86,
  output         OPIN_87,
  output         OPIN_88,
  input          clock,
  input          reset,
  input  [193:0] configBits,
  input          loopBreak,
  input          gndLBouts
);
  wire  alu_clock; // @[CLBlut4N10Mul.scala 45:53]
  wire  alu_reset; // @[CLBlut4N10Mul.scala 45:53]
  wire [15:0] alu_io_i0; // @[CLBlut4N10Mul.scala 45:53]
  wire [15:0] alu_io_i1; // @[CLBlut4N10Mul.scala 45:53]
  wire [31:0] alu_io_ib32; // @[CLBlut4N10Mul.scala 45:53]
  wire [7:0] alu_io_ctrl; // @[CLBlut4N10Mul.scala 45:53]
  wire [15:0] alu_io_q; // @[CLBlut4N10Mul.scala 45:53]
  wire [31:0] alu_io_config; // @[CLBlut4N10Mul.scala 45:53]
  wire  alu_io_gndOuts; // @[CLBlut4N10Mul.scala 45:53]
  wire  alu_io_clkEnb; // @[CLBlut4N10Mul.scala 45:53]
  wire  alu_io_loopBreak; // @[CLBlut4N10Mul.scala 45:53]
  wire  BLE_0_clock; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_0_reset; // @[CLBlut4N10Mul.scala 65:48]
  wire [19:0] BLE_0_io_config; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_0_io_in_0; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_0_io_in_1; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_0_io_in_2; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_0_io_in_3; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_0_io_outR; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_0_io_outT; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_0_io_gndOuts; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_0_io_clkEnb; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_0_io_loopBreak; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_clock; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_reset; // @[CLBlut4N10Mul.scala 65:48]
  wire [19:0] BLE_1_io_config; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_io_in_0; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_io_in_1; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_io_in_2; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_io_in_3; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_io_outR; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_io_outT; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_io_gndOuts; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_io_clkEnb; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_1_io_loopBreak; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_clock; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_reset; // @[CLBlut4N10Mul.scala 65:48]
  wire [19:0] BLE_2_io_config; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_io_in_0; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_io_in_1; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_io_in_2; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_io_in_3; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_io_outR; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_io_outT; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_io_gndOuts; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_io_clkEnb; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_2_io_loopBreak; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_clock; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_reset; // @[CLBlut4N10Mul.scala 65:48]
  wire [19:0] BLE_3_io_config; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_io_in_0; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_io_in_1; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_io_in_2; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_io_in_3; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_io_outR; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_io_outT; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_io_gndOuts; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_io_clkEnb; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_3_io_loopBreak; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_clock; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_reset; // @[CLBlut4N10Mul.scala 65:48]
  wire [19:0] BLE_4_io_config; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_io_in_0; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_io_in_1; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_io_in_2; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_io_in_3; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_io_outR; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_io_outT; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_io_gndOuts; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_io_clkEnb; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_4_io_loopBreak; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_clock; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_reset; // @[CLBlut4N10Mul.scala 65:48]
  wire [19:0] BLE_5_io_config; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_io_in_0; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_io_in_1; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_io_in_2; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_io_in_3; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_io_outR; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_io_outT; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_io_gndOuts; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_io_clkEnb; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_5_io_loopBreak; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_clock; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_reset; // @[CLBlut4N10Mul.scala 65:48]
  wire [19:0] BLE_6_io_config; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_io_in_0; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_io_in_1; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_io_in_2; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_io_in_3; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_io_outR; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_io_outT; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_io_gndOuts; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_io_clkEnb; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_6_io_loopBreak; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_clock; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_reset; // @[CLBlut4N10Mul.scala 65:48]
  wire [19:0] BLE_7_io_config; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_io_in_0; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_io_in_1; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_io_in_2; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_io_in_3; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_io_outR; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_io_outT; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_io_gndOuts; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_io_clkEnb; // @[CLBlut4N10Mul.scala 65:48]
  wire  BLE_7_io_loopBreak; // @[CLBlut4N10Mul.scala 65:48]
  wire [7:0] I_0 = {IPIN_7,IPIN_6,IPIN_5,IPIN_4,IPIN_3,IPIN_2,IPIN_1,IPIN_0}; // @[CLBlut4N10Mul.scala 35:92]
  wire [7:0] I_1 = {IPIN_15,IPIN_14,IPIN_13,IPIN_12,IPIN_11,IPIN_10,IPIN_9,IPIN_8}; // @[CLBlut4N10Mul.scala 35:92]
  wire [7:0] I_2 = {IPIN_23,IPIN_22,IPIN_21,IPIN_20,IPIN_19,IPIN_18,IPIN_17,IPIN_16}; // @[CLBlut4N10Mul.scala 35:92]
  wire [7:0] I_3 = {IPIN_31,IPIN_30,IPIN_29,IPIN_28,IPIN_27,IPIN_26,IPIN_25,IPIN_24}; // @[CLBlut4N10Mul.scala 35:92]
  wire  OAlu_0 = alu_io_q[0]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_0 = BLE_0_io_outR; // @[CLBlut4N10Mul.scala 38:18 70:15]
  wire  OAlu_1 = alu_io_q[1]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_1 = BLE_1_io_outR; // @[CLBlut4N10Mul.scala 38:18 70:15]
  wire  OAlu_2 = alu_io_q[2]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_2 = BLE_2_io_outR; // @[CLBlut4N10Mul.scala 38:18 70:15]
  wire  OAlu_3 = alu_io_q[3]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_3 = BLE_3_io_outR; // @[CLBlut4N10Mul.scala 38:18 70:15]
  wire  OAlu_4 = alu_io_q[4]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_4 = BLE_4_io_outR; // @[CLBlut4N10Mul.scala 38:18 70:15]
  wire  OAlu_5 = alu_io_q[5]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_5 = BLE_5_io_outR; // @[CLBlut4N10Mul.scala 38:18 70:15]
  wire  OAlu_6 = alu_io_q[6]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_6 = BLE_6_io_outR; // @[CLBlut4N10Mul.scala 38:18 70:15]
  wire  OAlu_7 = alu_io_q[7]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_7 = BLE_7_io_outR; // @[CLBlut4N10Mul.scala 38:18 70:15]
  wire  OAlu_8 = alu_io_q[8]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_8 = BLE_0_io_outT; // @[CLBlut4N10Mul.scala 38:18 71:17]
  wire  OAlu_9 = alu_io_q[9]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_9 = BLE_1_io_outT; // @[CLBlut4N10Mul.scala 38:18 71:17]
  wire  OAlu_10 = alu_io_q[10]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_10 = BLE_2_io_outT; // @[CLBlut4N10Mul.scala 38:18 71:17]
  wire  OAlu_11 = alu_io_q[11]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_11 = BLE_3_io_outT; // @[CLBlut4N10Mul.scala 38:18 71:17]
  wire  OAlu_12 = alu_io_q[12]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_12 = BLE_4_io_outT; // @[CLBlut4N10Mul.scala 38:18 71:17]
  wire  OAlu_13 = alu_io_q[13]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_13 = BLE_5_io_outT; // @[CLBlut4N10Mul.scala 38:18 71:17]
  wire  OAlu_14 = alu_io_q[14]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_14 = BLE_6_io_outT; // @[CLBlut4N10Mul.scala 38:18 71:17]
  wire  OAlu_15 = alu_io_q[15]; // @[CLBlut4N10Mul.scala 51:50]
  wire  OClb_15 = BLE_7_io_outT; // @[CLBlut4N10Mul.scala 38:18 71:17]
  wire [8:0] IPINsasUint_lo_lo_lo = {IPIN_8,IPIN_7,IPIN_6,IPIN_5,IPIN_4,IPIN_3,IPIN_2,IPIN_1,IPIN_0}; // @[CLBlut4N10Mul.scala 44:50]
  wire [17:0] IPINsasUint_lo_lo = {IPIN_17,IPIN_16,IPIN_15,IPIN_14,IPIN_13,IPIN_12,IPIN_11,IPIN_10,IPIN_9,
    IPINsasUint_lo_lo_lo}; // @[CLBlut4N10Mul.scala 44:50]
  wire [8:0] IPINsasUint_lo_hi_lo = {IPIN_26,IPIN_25,IPIN_24,IPIN_23,IPIN_22,IPIN_21,IPIN_20,IPIN_19,IPIN_18}; // @[CLBlut4N10Mul.scala 44:50]
  wire [17:0] IPINsasUint_lo_hi = {IPIN_35,IPIN_34,IPIN_33,IPIN_32,IPIN_31,IPIN_30,IPIN_29,IPIN_28,IPIN_27,
    IPINsasUint_lo_hi_lo}; // @[CLBlut4N10Mul.scala 44:50]
  wire [8:0] IPINsasUint_hi_lo_lo = {IPIN_44,IPIN_43,IPIN_42,IPIN_41,IPIN_40,IPIN_39,IPIN_38,IPIN_37,IPIN_36}; // @[CLBlut4N10Mul.scala 44:50]
  wire [17:0] IPINsasUint_hi_lo = {IPIN_53,IPIN_52,IPIN_51,IPIN_50,IPIN_49,IPIN_48,IPIN_47,IPIN_46,IPIN_45,
    IPINsasUint_hi_lo_lo}; // @[CLBlut4N10Mul.scala 44:50]
  wire [8:0] IPINsasUint_hi_hi_lo = {IPIN_62,IPIN_61,IPIN_60,IPIN_59,IPIN_58,IPIN_57,IPIN_56,IPIN_55,IPIN_54}; // @[CLBlut4N10Mul.scala 44:50]
  wire [17:0] IPINsasUint_hi_hi = {IPIN_71,IPIN_70,IPIN_69,IPIN_68,IPIN_67,IPIN_66,IPIN_65,IPIN_64,IPIN_63,
    IPINsasUint_hi_hi_lo}; // @[CLBlut4N10Mul.scala 44:50]
  wire [71:0] IPINsasUint = {IPINsasUint_hi_hi,IPINsasUint_hi_lo,IPINsasUint_lo_hi,IPINsasUint_lo_lo}; // @[CLBlut4N10Mul.scala 44:50]
  wire [1:0] _BLE_0_io_in_0_T_2 = {configBits[19],configBits[18]}; // @[Cat.scala 31:58]
  wire  _BLE_0_io_in_0_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_0[2] : I_0[2]; // @[Mux.scala 81:58]
  wire  _BLE_0_io_in_0_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_0[1] : _BLE_0_io_in_0_T_8; // @[Mux.scala 81:58]
  wire  _BLE_0_io_in_1_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_1[2] : I_1[2]; // @[Mux.scala 81:58]
  wire  _BLE_0_io_in_1_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_1[1] : _BLE_0_io_in_1_T_8; // @[Mux.scala 81:58]
  wire  _BLE_0_io_in_2_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_2[2] : I_2[2]; // @[Mux.scala 81:58]
  wire  _BLE_0_io_in_2_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_2[1] : _BLE_0_io_in_2_T_8; // @[Mux.scala 81:58]
  wire  _BLE_0_io_in_3_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_3[2] : I_3[2]; // @[Mux.scala 81:58]
  wire  _BLE_0_io_in_3_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_3[1] : _BLE_0_io_in_3_T_8; // @[Mux.scala 81:58]
  wire  _BLE_1_io_in_0_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_0[3] : I_0[3]; // @[Mux.scala 81:58]
  wire  _BLE_1_io_in_0_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_0[2] : _BLE_1_io_in_0_T_8; // @[Mux.scala 81:58]
  wire  _BLE_1_io_in_1_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_1[3] : I_1[3]; // @[Mux.scala 81:58]
  wire  _BLE_1_io_in_1_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_1[2] : _BLE_1_io_in_1_T_8; // @[Mux.scala 81:58]
  wire  _BLE_1_io_in_2_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_2[3] : I_2[3]; // @[Mux.scala 81:58]
  wire  _BLE_1_io_in_2_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_2[2] : _BLE_1_io_in_2_T_8; // @[Mux.scala 81:58]
  wire  _BLE_1_io_in_3_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_3[3] : I_3[3]; // @[Mux.scala 81:58]
  wire  _BLE_1_io_in_3_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_3[2] : _BLE_1_io_in_3_T_8; // @[Mux.scala 81:58]
  wire  _BLE_2_io_in_0_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_0[4] : I_0[4]; // @[Mux.scala 81:58]
  wire  _BLE_2_io_in_0_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_0[3] : _BLE_2_io_in_0_T_8; // @[Mux.scala 81:58]
  wire  _BLE_2_io_in_1_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_1[4] : I_1[4]; // @[Mux.scala 81:58]
  wire  _BLE_2_io_in_1_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_1[3] : _BLE_2_io_in_1_T_8; // @[Mux.scala 81:58]
  wire  _BLE_2_io_in_2_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_2[4] : I_2[4]; // @[Mux.scala 81:58]
  wire  _BLE_2_io_in_2_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_2[3] : _BLE_2_io_in_2_T_8; // @[Mux.scala 81:58]
  wire  _BLE_2_io_in_3_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_3[4] : I_3[4]; // @[Mux.scala 81:58]
  wire  _BLE_2_io_in_3_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_3[3] : _BLE_2_io_in_3_T_8; // @[Mux.scala 81:58]
  wire  _BLE_3_io_in_0_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_0[5] : I_0[5]; // @[Mux.scala 81:58]
  wire  _BLE_3_io_in_0_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_0[4] : _BLE_3_io_in_0_T_8; // @[Mux.scala 81:58]
  wire  _BLE_3_io_in_1_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_1[5] : I_1[5]; // @[Mux.scala 81:58]
  wire  _BLE_3_io_in_1_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_1[4] : _BLE_3_io_in_1_T_8; // @[Mux.scala 81:58]
  wire  _BLE_3_io_in_2_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_2[5] : I_2[5]; // @[Mux.scala 81:58]
  wire  _BLE_3_io_in_2_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_2[4] : _BLE_3_io_in_2_T_8; // @[Mux.scala 81:58]
  wire  _BLE_3_io_in_3_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_3[5] : I_3[5]; // @[Mux.scala 81:58]
  wire  _BLE_3_io_in_3_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_3[4] : _BLE_3_io_in_3_T_8; // @[Mux.scala 81:58]
  wire  _BLE_4_io_in_0_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_0[6] : I_0[6]; // @[Mux.scala 81:58]
  wire  _BLE_4_io_in_0_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_0[5] : _BLE_4_io_in_0_T_8; // @[Mux.scala 81:58]
  wire  _BLE_4_io_in_1_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_1[6] : I_1[6]; // @[Mux.scala 81:58]
  wire  _BLE_4_io_in_1_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_1[5] : _BLE_4_io_in_1_T_8; // @[Mux.scala 81:58]
  wire  _BLE_4_io_in_2_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_2[6] : I_2[6]; // @[Mux.scala 81:58]
  wire  _BLE_4_io_in_2_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_2[5] : _BLE_4_io_in_2_T_8; // @[Mux.scala 81:58]
  wire  _BLE_4_io_in_3_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_3[6] : I_3[6]; // @[Mux.scala 81:58]
  wire  _BLE_4_io_in_3_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_3[5] : _BLE_4_io_in_3_T_8; // @[Mux.scala 81:58]
  wire  _BLE_5_io_in_0_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_0[7] : I_0[7]; // @[Mux.scala 81:58]
  wire  _BLE_5_io_in_0_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_0[6] : _BLE_5_io_in_0_T_8; // @[Mux.scala 81:58]
  wire  _BLE_5_io_in_1_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_1[7] : I_1[7]; // @[Mux.scala 81:58]
  wire  _BLE_5_io_in_1_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_1[6] : _BLE_5_io_in_1_T_8; // @[Mux.scala 81:58]
  wire  _BLE_5_io_in_2_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_2[7] : I_2[7]; // @[Mux.scala 81:58]
  wire  _BLE_5_io_in_2_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_2[6] : _BLE_5_io_in_2_T_8; // @[Mux.scala 81:58]
  wire  _BLE_5_io_in_3_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_3[7] : I_3[7]; // @[Mux.scala 81:58]
  wire  _BLE_5_io_in_3_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_3[6] : _BLE_5_io_in_3_T_8; // @[Mux.scala 81:58]
  wire  _BLE_6_io_in_0_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_0[0] : I_0[0]; // @[Mux.scala 81:58]
  wire  _BLE_6_io_in_0_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_0[7] : _BLE_6_io_in_0_T_8; // @[Mux.scala 81:58]
  wire  _BLE_6_io_in_1_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_1[0] : I_1[0]; // @[Mux.scala 81:58]
  wire  _BLE_6_io_in_1_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_1[7] : _BLE_6_io_in_1_T_8; // @[Mux.scala 81:58]
  wire  _BLE_6_io_in_2_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_2[0] : I_2[0]; // @[Mux.scala 81:58]
  wire  _BLE_6_io_in_2_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_2[7] : _BLE_6_io_in_2_T_8; // @[Mux.scala 81:58]
  wire  _BLE_6_io_in_3_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_3[0] : I_3[0]; // @[Mux.scala 81:58]
  wire  _BLE_6_io_in_3_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_3[7] : _BLE_6_io_in_3_T_8; // @[Mux.scala 81:58]
  wire  _BLE_7_io_in_0_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_0[1] : I_0[1]; // @[Mux.scala 81:58]
  wire  _BLE_7_io_in_0_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_0[0] : _BLE_7_io_in_0_T_8; // @[Mux.scala 81:58]
  wire  _BLE_7_io_in_1_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_1[1] : I_1[1]; // @[Mux.scala 81:58]
  wire  _BLE_7_io_in_1_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_1[0] : _BLE_7_io_in_1_T_8; // @[Mux.scala 81:58]
  wire  _BLE_7_io_in_2_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_2[1] : I_2[1]; // @[Mux.scala 81:58]
  wire  _BLE_7_io_in_2_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_2[0] : _BLE_7_io_in_2_T_8; // @[Mux.scala 81:58]
  wire  _BLE_7_io_in_3_T_8 = 2'h2 == _BLE_0_io_in_0_T_2 ? I_3[1] : I_3[1]; // @[Mux.scala 81:58]
  wire  _BLE_7_io_in_3_T_10 = 2'h1 == _BLE_0_io_in_0_T_2 ? I_3[0] : _BLE_7_io_in_3_T_8; // @[Mux.scala 81:58]
  AluMul alu ( // @[CLBlut4N10Mul.scala 45:53]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_i0(alu_io_i0),
    .io_i1(alu_io_i1),
    .io_ib32(alu_io_ib32),
    .io_ctrl(alu_io_ctrl),
    .io_q(alu_io_q),
    .io_config(alu_io_config),
    .io_gndOuts(alu_io_gndOuts),
    .io_clkEnb(alu_io_clkEnb),
    .io_loopBreak(alu_io_loopBreak)
  );
  Ble4 BLE_0 ( // @[CLBlut4N10Mul.scala 65:48]
    .clock(BLE_0_clock),
    .reset(BLE_0_reset),
    .io_config(BLE_0_io_config),
    .io_in_0(BLE_0_io_in_0),
    .io_in_1(BLE_0_io_in_1),
    .io_in_2(BLE_0_io_in_2),
    .io_in_3(BLE_0_io_in_3),
    .io_outR(BLE_0_io_outR),
    .io_outT(BLE_0_io_outT),
    .io_gndOuts(BLE_0_io_gndOuts),
    .io_clkEnb(BLE_0_io_clkEnb),
    .io_loopBreak(BLE_0_io_loopBreak)
  );
  Ble4 BLE_1 ( // @[CLBlut4N10Mul.scala 65:48]
    .clock(BLE_1_clock),
    .reset(BLE_1_reset),
    .io_config(BLE_1_io_config),
    .io_in_0(BLE_1_io_in_0),
    .io_in_1(BLE_1_io_in_1),
    .io_in_2(BLE_1_io_in_2),
    .io_in_3(BLE_1_io_in_3),
    .io_outR(BLE_1_io_outR),
    .io_outT(BLE_1_io_outT),
    .io_gndOuts(BLE_1_io_gndOuts),
    .io_clkEnb(BLE_1_io_clkEnb),
    .io_loopBreak(BLE_1_io_loopBreak)
  );
  Ble4 BLE_2 ( // @[CLBlut4N10Mul.scala 65:48]
    .clock(BLE_2_clock),
    .reset(BLE_2_reset),
    .io_config(BLE_2_io_config),
    .io_in_0(BLE_2_io_in_0),
    .io_in_1(BLE_2_io_in_1),
    .io_in_2(BLE_2_io_in_2),
    .io_in_3(BLE_2_io_in_3),
    .io_outR(BLE_2_io_outR),
    .io_outT(BLE_2_io_outT),
    .io_gndOuts(BLE_2_io_gndOuts),
    .io_clkEnb(BLE_2_io_clkEnb),
    .io_loopBreak(BLE_2_io_loopBreak)
  );
  Ble4 BLE_3 ( // @[CLBlut4N10Mul.scala 65:48]
    .clock(BLE_3_clock),
    .reset(BLE_3_reset),
    .io_config(BLE_3_io_config),
    .io_in_0(BLE_3_io_in_0),
    .io_in_1(BLE_3_io_in_1),
    .io_in_2(BLE_3_io_in_2),
    .io_in_3(BLE_3_io_in_3),
    .io_outR(BLE_3_io_outR),
    .io_outT(BLE_3_io_outT),
    .io_gndOuts(BLE_3_io_gndOuts),
    .io_clkEnb(BLE_3_io_clkEnb),
    .io_loopBreak(BLE_3_io_loopBreak)
  );
  Ble4 BLE_4 ( // @[CLBlut4N10Mul.scala 65:48]
    .clock(BLE_4_clock),
    .reset(BLE_4_reset),
    .io_config(BLE_4_io_config),
    .io_in_0(BLE_4_io_in_0),
    .io_in_1(BLE_4_io_in_1),
    .io_in_2(BLE_4_io_in_2),
    .io_in_3(BLE_4_io_in_3),
    .io_outR(BLE_4_io_outR),
    .io_outT(BLE_4_io_outT),
    .io_gndOuts(BLE_4_io_gndOuts),
    .io_clkEnb(BLE_4_io_clkEnb),
    .io_loopBreak(BLE_4_io_loopBreak)
  );
  Ble4 BLE_5 ( // @[CLBlut4N10Mul.scala 65:48]
    .clock(BLE_5_clock),
    .reset(BLE_5_reset),
    .io_config(BLE_5_io_config),
    .io_in_0(BLE_5_io_in_0),
    .io_in_1(BLE_5_io_in_1),
    .io_in_2(BLE_5_io_in_2),
    .io_in_3(BLE_5_io_in_3),
    .io_outR(BLE_5_io_outR),
    .io_outT(BLE_5_io_outT),
    .io_gndOuts(BLE_5_io_gndOuts),
    .io_clkEnb(BLE_5_io_clkEnb),
    .io_loopBreak(BLE_5_io_loopBreak)
  );
  Ble4 BLE_6 ( // @[CLBlut4N10Mul.scala 65:48]
    .clock(BLE_6_clock),
    .reset(BLE_6_reset),
    .io_config(BLE_6_io_config),
    .io_in_0(BLE_6_io_in_0),
    .io_in_1(BLE_6_io_in_1),
    .io_in_2(BLE_6_io_in_2),
    .io_in_3(BLE_6_io_in_3),
    .io_outR(BLE_6_io_outR),
    .io_outT(BLE_6_io_outT),
    .io_gndOuts(BLE_6_io_gndOuts),
    .io_clkEnb(BLE_6_io_clkEnb),
    .io_loopBreak(BLE_6_io_loopBreak)
  );
  Ble4 BLE_7 ( // @[CLBlut4N10Mul.scala 65:48]
    .clock(BLE_7_clock),
    .reset(BLE_7_reset),
    .io_config(BLE_7_io_config),
    .io_in_0(BLE_7_io_in_0),
    .io_in_1(BLE_7_io_in_1),
    .io_in_2(BLE_7_io_in_2),
    .io_in_3(BLE_7_io_in_3),
    .io_outR(BLE_7_io_outR),
    .io_outT(BLE_7_io_outT),
    .io_gndOuts(BLE_7_io_gndOuts),
    .io_clkEnb(BLE_7_io_clkEnb),
    .io_loopBreak(BLE_7_io_loopBreak)
  );
  assign OPIN_73 = configBits[192] ? OAlu_0 & ~gndLBouts : OClb_0; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_74 = configBits[192] ? OAlu_1 & ~gndLBouts : OClb_1; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_75 = configBits[192] ? OAlu_2 & ~gndLBouts : OClb_2; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_76 = configBits[192] ? OAlu_3 & ~gndLBouts : OClb_3; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_77 = configBits[192] ? OAlu_4 & ~gndLBouts : OClb_4; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_78 = configBits[192] ? OAlu_5 & ~gndLBouts : OClb_5; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_79 = configBits[192] ? OAlu_6 & ~gndLBouts : OClb_6; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_80 = configBits[192] ? OAlu_7 & ~gndLBouts : OClb_7; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_81 = configBits[192] ? OAlu_8 & ~gndLBouts : OClb_8; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_82 = configBits[192] ? OAlu_9 & ~gndLBouts : OClb_9; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_83 = configBits[192] ? OAlu_10 & ~gndLBouts : OClb_10; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_84 = configBits[192] ? OAlu_11 & ~gndLBouts : OClb_11; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_85 = configBits[192] ? OAlu_12 & ~gndLBouts : OClb_12; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_86 = configBits[192] ? OAlu_13 & ~gndLBouts : OClb_13; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_87 = configBits[192] ? OAlu_14 & ~gndLBouts : OClb_14; // @[CLBlut4N10Mul.scala 40:15]
  assign OPIN_88 = configBits[192] ? OAlu_15 & ~gndLBouts : OClb_15; // @[CLBlut4N10Mul.scala 40:15]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_i0 = IPINsasUint[15:0]; // @[CLBlut4N10Mul.scala 47:27]
  assign alu_io_i1 = IPINsasUint[31:16]; // @[CLBlut4N10Mul.scala 48:27]
  assign alu_io_ib32 = IPINsasUint[71:40]; // @[CLBlut4N10Mul.scala 50:29]
  assign alu_io_ctrl = IPINsasUint[39:32]; // @[CLBlut4N10Mul.scala 49:29]
  assign alu_io_config = configBits[33:2]; // @[CLBlut4N10Mul.scala 55:30]
  assign alu_io_gndOuts = gndLBouts; // @[CLBlut4N10Mul.scala 54:18]
  assign alu_io_clkEnb = configBits[193]; // @[CLBlut4N10Mul.scala 53:30]
  assign alu_io_loopBreak = loopBreak; // @[CLBlut4N10Mul.scala 46:20]
  assign BLE_0_clock = clock;
  assign BLE_0_reset = reset;
  assign BLE_0_io_config = configBits[19:0]; // @[CLBlut4N10Mul.scala 67:38]
  assign BLE_0_io_in_0 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_0[0] : _BLE_0_io_in_0_T_10; // @[Mux.scala 81:58]
  assign BLE_0_io_in_1 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_1[0] : _BLE_0_io_in_1_T_10; // @[Mux.scala 81:58]
  assign BLE_0_io_in_2 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_2[0] : _BLE_0_io_in_2_T_10; // @[Mux.scala 81:58]
  assign BLE_0_io_in_3 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_3[0] : _BLE_0_io_in_3_T_10; // @[Mux.scala 81:58]
  assign BLE_0_io_gndOuts = gndLBouts; // @[CLBlut4N10Mul.scala 72:26]
  assign BLE_0_io_clkEnb = configBits[193]; // @[CLBlut4N10Mul.scala 73:38]
  assign BLE_0_io_loopBreak = loopBreak; // @[CLBlut4N10Mul.scala 74:28]
  assign BLE_1_clock = clock;
  assign BLE_1_reset = reset;
  assign BLE_1_io_config = configBits[39:20]; // @[CLBlut4N10Mul.scala 67:38]
  assign BLE_1_io_in_0 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_0[1] : _BLE_1_io_in_0_T_10; // @[Mux.scala 81:58]
  assign BLE_1_io_in_1 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_1[1] : _BLE_1_io_in_1_T_10; // @[Mux.scala 81:58]
  assign BLE_1_io_in_2 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_2[1] : _BLE_1_io_in_2_T_10; // @[Mux.scala 81:58]
  assign BLE_1_io_in_3 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_3[1] : _BLE_1_io_in_3_T_10; // @[Mux.scala 81:58]
  assign BLE_1_io_gndOuts = gndLBouts; // @[CLBlut4N10Mul.scala 72:26]
  assign BLE_1_io_clkEnb = configBits[193]; // @[CLBlut4N10Mul.scala 73:38]
  assign BLE_1_io_loopBreak = loopBreak; // @[CLBlut4N10Mul.scala 74:28]
  assign BLE_2_clock = clock;
  assign BLE_2_reset = reset;
  assign BLE_2_io_config = configBits[59:40]; // @[CLBlut4N10Mul.scala 67:38]
  assign BLE_2_io_in_0 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_0[2] : _BLE_2_io_in_0_T_10; // @[Mux.scala 81:58]
  assign BLE_2_io_in_1 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_1[2] : _BLE_2_io_in_1_T_10; // @[Mux.scala 81:58]
  assign BLE_2_io_in_2 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_2[2] : _BLE_2_io_in_2_T_10; // @[Mux.scala 81:58]
  assign BLE_2_io_in_3 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_3[2] : _BLE_2_io_in_3_T_10; // @[Mux.scala 81:58]
  assign BLE_2_io_gndOuts = gndLBouts; // @[CLBlut4N10Mul.scala 72:26]
  assign BLE_2_io_clkEnb = configBits[193]; // @[CLBlut4N10Mul.scala 73:38]
  assign BLE_2_io_loopBreak = loopBreak; // @[CLBlut4N10Mul.scala 74:28]
  assign BLE_3_clock = clock;
  assign BLE_3_reset = reset;
  assign BLE_3_io_config = configBits[79:60]; // @[CLBlut4N10Mul.scala 67:38]
  assign BLE_3_io_in_0 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_0[3] : _BLE_3_io_in_0_T_10; // @[Mux.scala 81:58]
  assign BLE_3_io_in_1 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_1[3] : _BLE_3_io_in_1_T_10; // @[Mux.scala 81:58]
  assign BLE_3_io_in_2 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_2[3] : _BLE_3_io_in_2_T_10; // @[Mux.scala 81:58]
  assign BLE_3_io_in_3 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_3[3] : _BLE_3_io_in_3_T_10; // @[Mux.scala 81:58]
  assign BLE_3_io_gndOuts = gndLBouts; // @[CLBlut4N10Mul.scala 72:26]
  assign BLE_3_io_clkEnb = configBits[193]; // @[CLBlut4N10Mul.scala 73:38]
  assign BLE_3_io_loopBreak = loopBreak; // @[CLBlut4N10Mul.scala 74:28]
  assign BLE_4_clock = clock;
  assign BLE_4_reset = reset;
  assign BLE_4_io_config = configBits[99:80]; // @[CLBlut4N10Mul.scala 67:38]
  assign BLE_4_io_in_0 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_0[4] : _BLE_4_io_in_0_T_10; // @[Mux.scala 81:58]
  assign BLE_4_io_in_1 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_1[4] : _BLE_4_io_in_1_T_10; // @[Mux.scala 81:58]
  assign BLE_4_io_in_2 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_2[4] : _BLE_4_io_in_2_T_10; // @[Mux.scala 81:58]
  assign BLE_4_io_in_3 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_3[4] : _BLE_4_io_in_3_T_10; // @[Mux.scala 81:58]
  assign BLE_4_io_gndOuts = gndLBouts; // @[CLBlut4N10Mul.scala 72:26]
  assign BLE_4_io_clkEnb = configBits[193]; // @[CLBlut4N10Mul.scala 73:38]
  assign BLE_4_io_loopBreak = loopBreak; // @[CLBlut4N10Mul.scala 74:28]
  assign BLE_5_clock = clock;
  assign BLE_5_reset = reset;
  assign BLE_5_io_config = configBits[119:100]; // @[CLBlut4N10Mul.scala 67:38]
  assign BLE_5_io_in_0 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_0[5] : _BLE_5_io_in_0_T_10; // @[Mux.scala 81:58]
  assign BLE_5_io_in_1 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_1[5] : _BLE_5_io_in_1_T_10; // @[Mux.scala 81:58]
  assign BLE_5_io_in_2 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_2[5] : _BLE_5_io_in_2_T_10; // @[Mux.scala 81:58]
  assign BLE_5_io_in_3 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_3[5] : _BLE_5_io_in_3_T_10; // @[Mux.scala 81:58]
  assign BLE_5_io_gndOuts = gndLBouts; // @[CLBlut4N10Mul.scala 72:26]
  assign BLE_5_io_clkEnb = configBits[193]; // @[CLBlut4N10Mul.scala 73:38]
  assign BLE_5_io_loopBreak = loopBreak; // @[CLBlut4N10Mul.scala 74:28]
  assign BLE_6_clock = clock;
  assign BLE_6_reset = reset;
  assign BLE_6_io_config = configBits[139:120]; // @[CLBlut4N10Mul.scala 67:38]
  assign BLE_6_io_in_0 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_0[6] : _BLE_6_io_in_0_T_10; // @[Mux.scala 81:58]
  assign BLE_6_io_in_1 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_1[6] : _BLE_6_io_in_1_T_10; // @[Mux.scala 81:58]
  assign BLE_6_io_in_2 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_2[6] : _BLE_6_io_in_2_T_10; // @[Mux.scala 81:58]
  assign BLE_6_io_in_3 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_3[6] : _BLE_6_io_in_3_T_10; // @[Mux.scala 81:58]
  assign BLE_6_io_gndOuts = gndLBouts; // @[CLBlut4N10Mul.scala 72:26]
  assign BLE_6_io_clkEnb = configBits[193]; // @[CLBlut4N10Mul.scala 73:38]
  assign BLE_6_io_loopBreak = loopBreak; // @[CLBlut4N10Mul.scala 74:28]
  assign BLE_7_clock = clock;
  assign BLE_7_reset = reset;
  assign BLE_7_io_config = configBits[159:140]; // @[CLBlut4N10Mul.scala 67:38]
  assign BLE_7_io_in_0 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_0[7] : _BLE_7_io_in_0_T_10; // @[Mux.scala 81:58]
  assign BLE_7_io_in_1 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_1[7] : _BLE_7_io_in_1_T_10; // @[Mux.scala 81:58]
  assign BLE_7_io_in_2 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_2[7] : _BLE_7_io_in_2_T_10; // @[Mux.scala 81:58]
  assign BLE_7_io_in_3 = 2'h0 == _BLE_0_io_in_0_T_2 ? I_3[7] : _BLE_7_io_in_3_T_10; // @[Mux.scala 81:58]
  assign BLE_7_io_gndOuts = gndLBouts; // @[CLBlut4N10Mul.scala 72:26]
  assign BLE_7_io_clkEnb = configBits[193]; // @[CLBlut4N10Mul.scala 73:38]
  assign BLE_7_io_loopBreak = loopBreak; // @[CLBlut4N10Mul.scala 74:28]
endmodule
module ScanConf_Tile_7_1_clbmultile(
  input          clock,
  output [655:0] ioBundle_confOut,
  input  [15:0]  ioBundle_scan_in,
  input          ioBundle_scan_en,
  output [15:0]  ioBundle_scan_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
`endif // RANDOMIZE_REG_INIT
  reg  confReg_0; // @[ScanConf.scala 32:20]
  reg  confReg_1; // @[ScanConf.scala 32:20]
  reg  confReg_2; // @[ScanConf.scala 32:20]
  reg  confReg_3; // @[ScanConf.scala 32:20]
  reg  confReg_4; // @[ScanConf.scala 32:20]
  reg  confReg_5; // @[ScanConf.scala 32:20]
  reg  confReg_6; // @[ScanConf.scala 32:20]
  reg  confReg_7; // @[ScanConf.scala 32:20]
  reg  confReg_8; // @[ScanConf.scala 32:20]
  reg  confReg_9; // @[ScanConf.scala 32:20]
  reg  confReg_10; // @[ScanConf.scala 32:20]
  reg  confReg_11; // @[ScanConf.scala 32:20]
  reg  confReg_12; // @[ScanConf.scala 32:20]
  reg  confReg_13; // @[ScanConf.scala 32:20]
  reg  confReg_14; // @[ScanConf.scala 32:20]
  reg  confReg_15; // @[ScanConf.scala 32:20]
  reg  confReg_16; // @[ScanConf.scala 32:20]
  reg  confReg_17; // @[ScanConf.scala 32:20]
  reg  confReg_18; // @[ScanConf.scala 32:20]
  reg  confReg_19; // @[ScanConf.scala 32:20]
  reg  confReg_20; // @[ScanConf.scala 32:20]
  reg  confReg_21; // @[ScanConf.scala 32:20]
  reg  confReg_22; // @[ScanConf.scala 32:20]
  reg  confReg_23; // @[ScanConf.scala 32:20]
  reg  confReg_24; // @[ScanConf.scala 32:20]
  reg  confReg_25; // @[ScanConf.scala 32:20]
  reg  confReg_26; // @[ScanConf.scala 32:20]
  reg  confReg_27; // @[ScanConf.scala 32:20]
  reg  confReg_28; // @[ScanConf.scala 32:20]
  reg  confReg_29; // @[ScanConf.scala 32:20]
  reg  confReg_30; // @[ScanConf.scala 32:20]
  reg  confReg_31; // @[ScanConf.scala 32:20]
  reg  confReg_32; // @[ScanConf.scala 32:20]
  reg  confReg_33; // @[ScanConf.scala 32:20]
  reg  confReg_34; // @[ScanConf.scala 32:20]
  reg  confReg_35; // @[ScanConf.scala 32:20]
  reg  confReg_36; // @[ScanConf.scala 32:20]
  reg  confReg_37; // @[ScanConf.scala 32:20]
  reg  confReg_38; // @[ScanConf.scala 32:20]
  reg  confReg_39; // @[ScanConf.scala 32:20]
  reg  confReg_40; // @[ScanConf.scala 32:20]
  reg  confReg_41; // @[ScanConf.scala 32:20]
  reg  confReg_42; // @[ScanConf.scala 32:20]
  reg  confReg_43; // @[ScanConf.scala 32:20]
  reg  confReg_44; // @[ScanConf.scala 32:20]
  reg  confReg_45; // @[ScanConf.scala 32:20]
  reg  confReg_46; // @[ScanConf.scala 32:20]
  reg  confReg_47; // @[ScanConf.scala 32:20]
  reg  confReg_48; // @[ScanConf.scala 32:20]
  reg  confReg_49; // @[ScanConf.scala 32:20]
  reg  confReg_50; // @[ScanConf.scala 32:20]
  reg  confReg_51; // @[ScanConf.scala 32:20]
  reg  confReg_52; // @[ScanConf.scala 32:20]
  reg  confReg_53; // @[ScanConf.scala 32:20]
  reg  confReg_54; // @[ScanConf.scala 32:20]
  reg  confReg_55; // @[ScanConf.scala 32:20]
  reg  confReg_56; // @[ScanConf.scala 32:20]
  reg  confReg_57; // @[ScanConf.scala 32:20]
  reg  confReg_58; // @[ScanConf.scala 32:20]
  reg  confReg_59; // @[ScanConf.scala 32:20]
  reg  confReg_60; // @[ScanConf.scala 32:20]
  reg  confReg_61; // @[ScanConf.scala 32:20]
  reg  confReg_62; // @[ScanConf.scala 32:20]
  reg  confReg_63; // @[ScanConf.scala 32:20]
  reg  confReg_64; // @[ScanConf.scala 32:20]
  reg  confReg_65; // @[ScanConf.scala 32:20]
  reg  confReg_66; // @[ScanConf.scala 32:20]
  reg  confReg_67; // @[ScanConf.scala 32:20]
  reg  confReg_68; // @[ScanConf.scala 32:20]
  reg  confReg_69; // @[ScanConf.scala 32:20]
  reg  confReg_70; // @[ScanConf.scala 32:20]
  reg  confReg_71; // @[ScanConf.scala 32:20]
  reg  confReg_72; // @[ScanConf.scala 32:20]
  reg  confReg_73; // @[ScanConf.scala 32:20]
  reg  confReg_74; // @[ScanConf.scala 32:20]
  reg  confReg_75; // @[ScanConf.scala 32:20]
  reg  confReg_76; // @[ScanConf.scala 32:20]
  reg  confReg_77; // @[ScanConf.scala 32:20]
  reg  confReg_78; // @[ScanConf.scala 32:20]
  reg  confReg_79; // @[ScanConf.scala 32:20]
  reg  confReg_80; // @[ScanConf.scala 32:20]
  reg  confReg_81; // @[ScanConf.scala 32:20]
  reg  confReg_82; // @[ScanConf.scala 32:20]
  reg  confReg_83; // @[ScanConf.scala 32:20]
  reg  confReg_84; // @[ScanConf.scala 32:20]
  reg  confReg_85; // @[ScanConf.scala 32:20]
  reg  confReg_86; // @[ScanConf.scala 32:20]
  reg  confReg_87; // @[ScanConf.scala 32:20]
  reg  confReg_88; // @[ScanConf.scala 32:20]
  reg  confReg_89; // @[ScanConf.scala 32:20]
  reg  confReg_90; // @[ScanConf.scala 32:20]
  reg  confReg_91; // @[ScanConf.scala 32:20]
  reg  confReg_92; // @[ScanConf.scala 32:20]
  reg  confReg_93; // @[ScanConf.scala 32:20]
  reg  confReg_94; // @[ScanConf.scala 32:20]
  reg  confReg_95; // @[ScanConf.scala 32:20]
  reg  confReg_96; // @[ScanConf.scala 32:20]
  reg  confReg_97; // @[ScanConf.scala 32:20]
  reg  confReg_98; // @[ScanConf.scala 32:20]
  reg  confReg_99; // @[ScanConf.scala 32:20]
  reg  confReg_100; // @[ScanConf.scala 32:20]
  reg  confReg_101; // @[ScanConf.scala 32:20]
  reg  confReg_102; // @[ScanConf.scala 32:20]
  reg  confReg_103; // @[ScanConf.scala 32:20]
  reg  confReg_104; // @[ScanConf.scala 32:20]
  reg  confReg_105; // @[ScanConf.scala 32:20]
  reg  confReg_106; // @[ScanConf.scala 32:20]
  reg  confReg_107; // @[ScanConf.scala 32:20]
  reg  confReg_108; // @[ScanConf.scala 32:20]
  reg  confReg_109; // @[ScanConf.scala 32:20]
  reg  confReg_110; // @[ScanConf.scala 32:20]
  reg  confReg_111; // @[ScanConf.scala 32:20]
  reg  confReg_112; // @[ScanConf.scala 32:20]
  reg  confReg_113; // @[ScanConf.scala 32:20]
  reg  confReg_114; // @[ScanConf.scala 32:20]
  reg  confReg_115; // @[ScanConf.scala 32:20]
  reg  confReg_116; // @[ScanConf.scala 32:20]
  reg  confReg_117; // @[ScanConf.scala 32:20]
  reg  confReg_118; // @[ScanConf.scala 32:20]
  reg  confReg_119; // @[ScanConf.scala 32:20]
  reg  confReg_120; // @[ScanConf.scala 32:20]
  reg  confReg_121; // @[ScanConf.scala 32:20]
  reg  confReg_122; // @[ScanConf.scala 32:20]
  reg  confReg_123; // @[ScanConf.scala 32:20]
  reg  confReg_124; // @[ScanConf.scala 32:20]
  reg  confReg_125; // @[ScanConf.scala 32:20]
  reg  confReg_126; // @[ScanConf.scala 32:20]
  reg  confReg_127; // @[ScanConf.scala 32:20]
  reg  confReg_128; // @[ScanConf.scala 32:20]
  reg  confReg_129; // @[ScanConf.scala 32:20]
  reg  confReg_130; // @[ScanConf.scala 32:20]
  reg  confReg_131; // @[ScanConf.scala 32:20]
  reg  confReg_132; // @[ScanConf.scala 32:20]
  reg  confReg_133; // @[ScanConf.scala 32:20]
  reg  confReg_134; // @[ScanConf.scala 32:20]
  reg  confReg_135; // @[ScanConf.scala 32:20]
  reg  confReg_136; // @[ScanConf.scala 32:20]
  reg  confReg_137; // @[ScanConf.scala 32:20]
  reg  confReg_138; // @[ScanConf.scala 32:20]
  reg  confReg_139; // @[ScanConf.scala 32:20]
  reg  confReg_140; // @[ScanConf.scala 32:20]
  reg  confReg_141; // @[ScanConf.scala 32:20]
  reg  confReg_142; // @[ScanConf.scala 32:20]
  reg  confReg_143; // @[ScanConf.scala 32:20]
  reg  confReg_144; // @[ScanConf.scala 32:20]
  reg  confReg_145; // @[ScanConf.scala 32:20]
  reg  confReg_146; // @[ScanConf.scala 32:20]
  reg  confReg_147; // @[ScanConf.scala 32:20]
  reg  confReg_148; // @[ScanConf.scala 32:20]
  reg  confReg_149; // @[ScanConf.scala 32:20]
  reg  confReg_150; // @[ScanConf.scala 32:20]
  reg  confReg_151; // @[ScanConf.scala 32:20]
  reg  confReg_152; // @[ScanConf.scala 32:20]
  reg  confReg_153; // @[ScanConf.scala 32:20]
  reg  confReg_154; // @[ScanConf.scala 32:20]
  reg  confReg_155; // @[ScanConf.scala 32:20]
  reg  confReg_156; // @[ScanConf.scala 32:20]
  reg  confReg_157; // @[ScanConf.scala 32:20]
  reg  confReg_158; // @[ScanConf.scala 32:20]
  reg  confReg_159; // @[ScanConf.scala 32:20]
  reg  confReg_160; // @[ScanConf.scala 32:20]
  reg  confReg_161; // @[ScanConf.scala 32:20]
  reg  confReg_162; // @[ScanConf.scala 32:20]
  reg  confReg_163; // @[ScanConf.scala 32:20]
  reg  confReg_164; // @[ScanConf.scala 32:20]
  reg  confReg_165; // @[ScanConf.scala 32:20]
  reg  confReg_166; // @[ScanConf.scala 32:20]
  reg  confReg_167; // @[ScanConf.scala 32:20]
  reg  confReg_168; // @[ScanConf.scala 32:20]
  reg  confReg_169; // @[ScanConf.scala 32:20]
  reg  confReg_170; // @[ScanConf.scala 32:20]
  reg  confReg_171; // @[ScanConf.scala 32:20]
  reg  confReg_172; // @[ScanConf.scala 32:20]
  reg  confReg_173; // @[ScanConf.scala 32:20]
  reg  confReg_174; // @[ScanConf.scala 32:20]
  reg  confReg_175; // @[ScanConf.scala 32:20]
  reg  confReg_176; // @[ScanConf.scala 32:20]
  reg  confReg_177; // @[ScanConf.scala 32:20]
  reg  confReg_178; // @[ScanConf.scala 32:20]
  reg  confReg_179; // @[ScanConf.scala 32:20]
  reg  confReg_180; // @[ScanConf.scala 32:20]
  reg  confReg_181; // @[ScanConf.scala 32:20]
  reg  confReg_182; // @[ScanConf.scala 32:20]
  reg  confReg_183; // @[ScanConf.scala 32:20]
  reg  confReg_184; // @[ScanConf.scala 32:20]
  reg  confReg_185; // @[ScanConf.scala 32:20]
  reg  confReg_186; // @[ScanConf.scala 32:20]
  reg  confReg_187; // @[ScanConf.scala 32:20]
  reg  confReg_188; // @[ScanConf.scala 32:20]
  reg  confReg_189; // @[ScanConf.scala 32:20]
  reg  confReg_190; // @[ScanConf.scala 32:20]
  reg  confReg_191; // @[ScanConf.scala 32:20]
  reg  confReg_192; // @[ScanConf.scala 32:20]
  reg  confReg_193; // @[ScanConf.scala 32:20]
  reg  confReg_194; // @[ScanConf.scala 32:20]
  reg  confReg_195; // @[ScanConf.scala 32:20]
  reg  confReg_196; // @[ScanConf.scala 32:20]
  reg  confReg_197; // @[ScanConf.scala 32:20]
  reg  confReg_198; // @[ScanConf.scala 32:20]
  reg  confReg_199; // @[ScanConf.scala 32:20]
  reg  confReg_200; // @[ScanConf.scala 32:20]
  reg  confReg_201; // @[ScanConf.scala 32:20]
  reg  confReg_202; // @[ScanConf.scala 32:20]
  reg  confReg_203; // @[ScanConf.scala 32:20]
  reg  confReg_204; // @[ScanConf.scala 32:20]
  reg  confReg_205; // @[ScanConf.scala 32:20]
  reg  confReg_206; // @[ScanConf.scala 32:20]
  reg  confReg_207; // @[ScanConf.scala 32:20]
  reg  confReg_208; // @[ScanConf.scala 32:20]
  reg  confReg_209; // @[ScanConf.scala 32:20]
  reg  confReg_210; // @[ScanConf.scala 32:20]
  reg  confReg_211; // @[ScanConf.scala 32:20]
  reg  confReg_212; // @[ScanConf.scala 32:20]
  reg  confReg_213; // @[ScanConf.scala 32:20]
  reg  confReg_214; // @[ScanConf.scala 32:20]
  reg  confReg_215; // @[ScanConf.scala 32:20]
  reg  confReg_216; // @[ScanConf.scala 32:20]
  reg  confReg_217; // @[ScanConf.scala 32:20]
  reg  confReg_218; // @[ScanConf.scala 32:20]
  reg  confReg_219; // @[ScanConf.scala 32:20]
  reg  confReg_220; // @[ScanConf.scala 32:20]
  reg  confReg_221; // @[ScanConf.scala 32:20]
  reg  confReg_222; // @[ScanConf.scala 32:20]
  reg  confReg_223; // @[ScanConf.scala 32:20]
  reg  confReg_224; // @[ScanConf.scala 32:20]
  reg  confReg_225; // @[ScanConf.scala 32:20]
  reg  confReg_226; // @[ScanConf.scala 32:20]
  reg  confReg_227; // @[ScanConf.scala 32:20]
  reg  confReg_228; // @[ScanConf.scala 32:20]
  reg  confReg_229; // @[ScanConf.scala 32:20]
  reg  confReg_230; // @[ScanConf.scala 32:20]
  reg  confReg_231; // @[ScanConf.scala 32:20]
  reg  confReg_232; // @[ScanConf.scala 32:20]
  reg  confReg_233; // @[ScanConf.scala 32:20]
  reg  confReg_234; // @[ScanConf.scala 32:20]
  reg  confReg_235; // @[ScanConf.scala 32:20]
  reg  confReg_236; // @[ScanConf.scala 32:20]
  reg  confReg_237; // @[ScanConf.scala 32:20]
  reg  confReg_238; // @[ScanConf.scala 32:20]
  reg  confReg_239; // @[ScanConf.scala 32:20]
  reg  confReg_240; // @[ScanConf.scala 32:20]
  reg  confReg_241; // @[ScanConf.scala 32:20]
  reg  confReg_242; // @[ScanConf.scala 32:20]
  reg  confReg_243; // @[ScanConf.scala 32:20]
  reg  confReg_244; // @[ScanConf.scala 32:20]
  reg  confReg_245; // @[ScanConf.scala 32:20]
  reg  confReg_246; // @[ScanConf.scala 32:20]
  reg  confReg_247; // @[ScanConf.scala 32:20]
  reg  confReg_248; // @[ScanConf.scala 32:20]
  reg  confReg_249; // @[ScanConf.scala 32:20]
  reg  confReg_250; // @[ScanConf.scala 32:20]
  reg  confReg_251; // @[ScanConf.scala 32:20]
  reg  confReg_252; // @[ScanConf.scala 32:20]
  reg  confReg_253; // @[ScanConf.scala 32:20]
  reg  confReg_254; // @[ScanConf.scala 32:20]
  reg  confReg_255; // @[ScanConf.scala 32:20]
  reg  confReg_256; // @[ScanConf.scala 32:20]
  reg  confReg_257; // @[ScanConf.scala 32:20]
  reg  confReg_258; // @[ScanConf.scala 32:20]
  reg  confReg_259; // @[ScanConf.scala 32:20]
  reg  confReg_260; // @[ScanConf.scala 32:20]
  reg  confReg_261; // @[ScanConf.scala 32:20]
  reg  confReg_262; // @[ScanConf.scala 32:20]
  reg  confReg_263; // @[ScanConf.scala 32:20]
  reg  confReg_264; // @[ScanConf.scala 32:20]
  reg  confReg_265; // @[ScanConf.scala 32:20]
  reg  confReg_266; // @[ScanConf.scala 32:20]
  reg  confReg_267; // @[ScanConf.scala 32:20]
  reg  confReg_268; // @[ScanConf.scala 32:20]
  reg  confReg_269; // @[ScanConf.scala 32:20]
  reg  confReg_270; // @[ScanConf.scala 32:20]
  reg  confReg_271; // @[ScanConf.scala 32:20]
  reg  confReg_272; // @[ScanConf.scala 32:20]
  reg  confReg_273; // @[ScanConf.scala 32:20]
  reg  confReg_274; // @[ScanConf.scala 32:20]
  reg  confReg_275; // @[ScanConf.scala 32:20]
  reg  confReg_276; // @[ScanConf.scala 32:20]
  reg  confReg_277; // @[ScanConf.scala 32:20]
  reg  confReg_278; // @[ScanConf.scala 32:20]
  reg  confReg_279; // @[ScanConf.scala 32:20]
  reg  confReg_280; // @[ScanConf.scala 32:20]
  reg  confReg_281; // @[ScanConf.scala 32:20]
  reg  confReg_282; // @[ScanConf.scala 32:20]
  reg  confReg_283; // @[ScanConf.scala 32:20]
  reg  confReg_284; // @[ScanConf.scala 32:20]
  reg  confReg_285; // @[ScanConf.scala 32:20]
  reg  confReg_286; // @[ScanConf.scala 32:20]
  reg  confReg_287; // @[ScanConf.scala 32:20]
  reg  confReg_288; // @[ScanConf.scala 32:20]
  reg  confReg_289; // @[ScanConf.scala 32:20]
  reg  confReg_290; // @[ScanConf.scala 32:20]
  reg  confReg_291; // @[ScanConf.scala 32:20]
  reg  confReg_292; // @[ScanConf.scala 32:20]
  reg  confReg_293; // @[ScanConf.scala 32:20]
  reg  confReg_294; // @[ScanConf.scala 32:20]
  reg  confReg_295; // @[ScanConf.scala 32:20]
  reg  confReg_296; // @[ScanConf.scala 32:20]
  reg  confReg_297; // @[ScanConf.scala 32:20]
  reg  confReg_298; // @[ScanConf.scala 32:20]
  reg  confReg_299; // @[ScanConf.scala 32:20]
  reg  confReg_300; // @[ScanConf.scala 32:20]
  reg  confReg_301; // @[ScanConf.scala 32:20]
  reg  confReg_302; // @[ScanConf.scala 32:20]
  reg  confReg_303; // @[ScanConf.scala 32:20]
  reg  confReg_304; // @[ScanConf.scala 32:20]
  reg  confReg_305; // @[ScanConf.scala 32:20]
  reg  confReg_306; // @[ScanConf.scala 32:20]
  reg  confReg_307; // @[ScanConf.scala 32:20]
  reg  confReg_308; // @[ScanConf.scala 32:20]
  reg  confReg_309; // @[ScanConf.scala 32:20]
  reg  confReg_310; // @[ScanConf.scala 32:20]
  reg  confReg_311; // @[ScanConf.scala 32:20]
  reg  confReg_312; // @[ScanConf.scala 32:20]
  reg  confReg_313; // @[ScanConf.scala 32:20]
  reg  confReg_314; // @[ScanConf.scala 32:20]
  reg  confReg_315; // @[ScanConf.scala 32:20]
  reg  confReg_316; // @[ScanConf.scala 32:20]
  reg  confReg_317; // @[ScanConf.scala 32:20]
  reg  confReg_318; // @[ScanConf.scala 32:20]
  reg  confReg_319; // @[ScanConf.scala 32:20]
  reg  confReg_320; // @[ScanConf.scala 32:20]
  reg  confReg_321; // @[ScanConf.scala 32:20]
  reg  confReg_322; // @[ScanConf.scala 32:20]
  reg  confReg_323; // @[ScanConf.scala 32:20]
  reg  confReg_324; // @[ScanConf.scala 32:20]
  reg  confReg_325; // @[ScanConf.scala 32:20]
  reg  confReg_326; // @[ScanConf.scala 32:20]
  reg  confReg_327; // @[ScanConf.scala 32:20]
  reg  confReg_328; // @[ScanConf.scala 32:20]
  reg  confReg_329; // @[ScanConf.scala 32:20]
  reg  confReg_330; // @[ScanConf.scala 32:20]
  reg  confReg_331; // @[ScanConf.scala 32:20]
  reg  confReg_332; // @[ScanConf.scala 32:20]
  reg  confReg_333; // @[ScanConf.scala 32:20]
  reg  confReg_334; // @[ScanConf.scala 32:20]
  reg  confReg_335; // @[ScanConf.scala 32:20]
  reg  confReg_336; // @[ScanConf.scala 32:20]
  reg  confReg_337; // @[ScanConf.scala 32:20]
  reg  confReg_338; // @[ScanConf.scala 32:20]
  reg  confReg_339; // @[ScanConf.scala 32:20]
  reg  confReg_340; // @[ScanConf.scala 32:20]
  reg  confReg_341; // @[ScanConf.scala 32:20]
  reg  confReg_342; // @[ScanConf.scala 32:20]
  reg  confReg_343; // @[ScanConf.scala 32:20]
  reg  confReg_344; // @[ScanConf.scala 32:20]
  reg  confReg_345; // @[ScanConf.scala 32:20]
  reg  confReg_346; // @[ScanConf.scala 32:20]
  reg  confReg_347; // @[ScanConf.scala 32:20]
  reg  confReg_348; // @[ScanConf.scala 32:20]
  reg  confReg_349; // @[ScanConf.scala 32:20]
  reg  confReg_350; // @[ScanConf.scala 32:20]
  reg  confReg_351; // @[ScanConf.scala 32:20]
  reg  confReg_352; // @[ScanConf.scala 32:20]
  reg  confReg_353; // @[ScanConf.scala 32:20]
  reg  confReg_354; // @[ScanConf.scala 32:20]
  reg  confReg_355; // @[ScanConf.scala 32:20]
  reg  confReg_356; // @[ScanConf.scala 32:20]
  reg  confReg_357; // @[ScanConf.scala 32:20]
  reg  confReg_358; // @[ScanConf.scala 32:20]
  reg  confReg_359; // @[ScanConf.scala 32:20]
  reg  confReg_360; // @[ScanConf.scala 32:20]
  reg  confReg_361; // @[ScanConf.scala 32:20]
  reg  confReg_362; // @[ScanConf.scala 32:20]
  reg  confReg_363; // @[ScanConf.scala 32:20]
  reg  confReg_364; // @[ScanConf.scala 32:20]
  reg  confReg_365; // @[ScanConf.scala 32:20]
  reg  confReg_366; // @[ScanConf.scala 32:20]
  reg  confReg_367; // @[ScanConf.scala 32:20]
  reg  confReg_368; // @[ScanConf.scala 32:20]
  reg  confReg_369; // @[ScanConf.scala 32:20]
  reg  confReg_370; // @[ScanConf.scala 32:20]
  reg  confReg_371; // @[ScanConf.scala 32:20]
  reg  confReg_372; // @[ScanConf.scala 32:20]
  reg  confReg_373; // @[ScanConf.scala 32:20]
  reg  confReg_374; // @[ScanConf.scala 32:20]
  reg  confReg_375; // @[ScanConf.scala 32:20]
  reg  confReg_376; // @[ScanConf.scala 32:20]
  reg  confReg_377; // @[ScanConf.scala 32:20]
  reg  confReg_378; // @[ScanConf.scala 32:20]
  reg  confReg_379; // @[ScanConf.scala 32:20]
  reg  confReg_380; // @[ScanConf.scala 32:20]
  reg  confReg_381; // @[ScanConf.scala 32:20]
  reg  confReg_382; // @[ScanConf.scala 32:20]
  reg  confReg_383; // @[ScanConf.scala 32:20]
  reg  confReg_384; // @[ScanConf.scala 32:20]
  reg  confReg_385; // @[ScanConf.scala 32:20]
  reg  confReg_386; // @[ScanConf.scala 32:20]
  reg  confReg_387; // @[ScanConf.scala 32:20]
  reg  confReg_388; // @[ScanConf.scala 32:20]
  reg  confReg_389; // @[ScanConf.scala 32:20]
  reg  confReg_390; // @[ScanConf.scala 32:20]
  reg  confReg_391; // @[ScanConf.scala 32:20]
  reg  confReg_392; // @[ScanConf.scala 32:20]
  reg  confReg_393; // @[ScanConf.scala 32:20]
  reg  confReg_394; // @[ScanConf.scala 32:20]
  reg  confReg_395; // @[ScanConf.scala 32:20]
  reg  confReg_396; // @[ScanConf.scala 32:20]
  reg  confReg_397; // @[ScanConf.scala 32:20]
  reg  confReg_398; // @[ScanConf.scala 32:20]
  reg  confReg_399; // @[ScanConf.scala 32:20]
  reg  confReg_400; // @[ScanConf.scala 32:20]
  reg  confReg_401; // @[ScanConf.scala 32:20]
  reg  confReg_402; // @[ScanConf.scala 32:20]
  reg  confReg_403; // @[ScanConf.scala 32:20]
  reg  confReg_404; // @[ScanConf.scala 32:20]
  reg  confReg_405; // @[ScanConf.scala 32:20]
  reg  confReg_406; // @[ScanConf.scala 32:20]
  reg  confReg_407; // @[ScanConf.scala 32:20]
  reg  confReg_408; // @[ScanConf.scala 32:20]
  reg  confReg_409; // @[ScanConf.scala 32:20]
  reg  confReg_410; // @[ScanConf.scala 32:20]
  reg  confReg_411; // @[ScanConf.scala 32:20]
  reg  confReg_412; // @[ScanConf.scala 32:20]
  reg  confReg_413; // @[ScanConf.scala 32:20]
  reg  confReg_414; // @[ScanConf.scala 32:20]
  reg  confReg_415; // @[ScanConf.scala 32:20]
  reg  confReg_416; // @[ScanConf.scala 32:20]
  reg  confReg_417; // @[ScanConf.scala 32:20]
  reg  confReg_418; // @[ScanConf.scala 32:20]
  reg  confReg_419; // @[ScanConf.scala 32:20]
  reg  confReg_420; // @[ScanConf.scala 32:20]
  reg  confReg_421; // @[ScanConf.scala 32:20]
  reg  confReg_422; // @[ScanConf.scala 32:20]
  reg  confReg_423; // @[ScanConf.scala 32:20]
  reg  confReg_424; // @[ScanConf.scala 32:20]
  reg  confReg_425; // @[ScanConf.scala 32:20]
  reg  confReg_426; // @[ScanConf.scala 32:20]
  reg  confReg_427; // @[ScanConf.scala 32:20]
  reg  confReg_428; // @[ScanConf.scala 32:20]
  reg  confReg_429; // @[ScanConf.scala 32:20]
  reg  confReg_430; // @[ScanConf.scala 32:20]
  reg  confReg_431; // @[ScanConf.scala 32:20]
  reg  confReg_432; // @[ScanConf.scala 32:20]
  reg  confReg_433; // @[ScanConf.scala 32:20]
  reg  confReg_434; // @[ScanConf.scala 32:20]
  reg  confReg_435; // @[ScanConf.scala 32:20]
  reg  confReg_436; // @[ScanConf.scala 32:20]
  reg  confReg_437; // @[ScanConf.scala 32:20]
  reg  confReg_438; // @[ScanConf.scala 32:20]
  reg  confReg_439; // @[ScanConf.scala 32:20]
  reg  confReg_440; // @[ScanConf.scala 32:20]
  reg  confReg_441; // @[ScanConf.scala 32:20]
  reg  confReg_442; // @[ScanConf.scala 32:20]
  reg  confReg_443; // @[ScanConf.scala 32:20]
  reg  confReg_444; // @[ScanConf.scala 32:20]
  reg  confReg_445; // @[ScanConf.scala 32:20]
  reg  confReg_446; // @[ScanConf.scala 32:20]
  reg  confReg_447; // @[ScanConf.scala 32:20]
  reg  confReg_448; // @[ScanConf.scala 32:20]
  reg  confReg_449; // @[ScanConf.scala 32:20]
  reg  confReg_450; // @[ScanConf.scala 32:20]
  reg  confReg_451; // @[ScanConf.scala 32:20]
  reg  confReg_452; // @[ScanConf.scala 32:20]
  reg  confReg_453; // @[ScanConf.scala 32:20]
  reg  confReg_454; // @[ScanConf.scala 32:20]
  reg  confReg_455; // @[ScanConf.scala 32:20]
  reg  confReg_456; // @[ScanConf.scala 32:20]
  reg  confReg_457; // @[ScanConf.scala 32:20]
  reg  confReg_458; // @[ScanConf.scala 32:20]
  reg  confReg_459; // @[ScanConf.scala 32:20]
  reg  confReg_460; // @[ScanConf.scala 32:20]
  reg  confReg_461; // @[ScanConf.scala 32:20]
  reg  confReg_462; // @[ScanConf.scala 32:20]
  reg  confReg_463; // @[ScanConf.scala 32:20]
  reg  confReg_464; // @[ScanConf.scala 32:20]
  reg  confReg_465; // @[ScanConf.scala 32:20]
  reg  confReg_466; // @[ScanConf.scala 32:20]
  reg  confReg_467; // @[ScanConf.scala 32:20]
  reg  confReg_468; // @[ScanConf.scala 32:20]
  reg  confReg_469; // @[ScanConf.scala 32:20]
  reg  confReg_470; // @[ScanConf.scala 32:20]
  reg  confReg_471; // @[ScanConf.scala 32:20]
  reg  confReg_472; // @[ScanConf.scala 32:20]
  reg  confReg_473; // @[ScanConf.scala 32:20]
  reg  confReg_474; // @[ScanConf.scala 32:20]
  reg  confReg_475; // @[ScanConf.scala 32:20]
  reg  confReg_476; // @[ScanConf.scala 32:20]
  reg  confReg_477; // @[ScanConf.scala 32:20]
  reg  confReg_478; // @[ScanConf.scala 32:20]
  reg  confReg_479; // @[ScanConf.scala 32:20]
  reg  confReg_480; // @[ScanConf.scala 32:20]
  reg  confReg_481; // @[ScanConf.scala 32:20]
  reg  confReg_482; // @[ScanConf.scala 32:20]
  reg  confReg_483; // @[ScanConf.scala 32:20]
  reg  confReg_484; // @[ScanConf.scala 32:20]
  reg  confReg_485; // @[ScanConf.scala 32:20]
  reg  confReg_486; // @[ScanConf.scala 32:20]
  reg  confReg_487; // @[ScanConf.scala 32:20]
  reg  confReg_488; // @[ScanConf.scala 32:20]
  reg  confReg_489; // @[ScanConf.scala 32:20]
  reg  confReg_490; // @[ScanConf.scala 32:20]
  reg  confReg_491; // @[ScanConf.scala 32:20]
  reg  confReg_492; // @[ScanConf.scala 32:20]
  reg  confReg_493; // @[ScanConf.scala 32:20]
  reg  confReg_494; // @[ScanConf.scala 32:20]
  reg  confReg_495; // @[ScanConf.scala 32:20]
  reg  confReg_496; // @[ScanConf.scala 32:20]
  reg  confReg_497; // @[ScanConf.scala 32:20]
  reg  confReg_498; // @[ScanConf.scala 32:20]
  reg  confReg_499; // @[ScanConf.scala 32:20]
  reg  confReg_500; // @[ScanConf.scala 32:20]
  reg  confReg_501; // @[ScanConf.scala 32:20]
  reg  confReg_502; // @[ScanConf.scala 32:20]
  reg  confReg_503; // @[ScanConf.scala 32:20]
  reg  confReg_504; // @[ScanConf.scala 32:20]
  reg  confReg_505; // @[ScanConf.scala 32:20]
  reg  confReg_506; // @[ScanConf.scala 32:20]
  reg  confReg_507; // @[ScanConf.scala 32:20]
  reg  confReg_508; // @[ScanConf.scala 32:20]
  reg  confReg_509; // @[ScanConf.scala 32:20]
  reg  confReg_510; // @[ScanConf.scala 32:20]
  reg  confReg_511; // @[ScanConf.scala 32:20]
  reg  confReg_512; // @[ScanConf.scala 32:20]
  reg  confReg_513; // @[ScanConf.scala 32:20]
  reg  confReg_514; // @[ScanConf.scala 32:20]
  reg  confReg_515; // @[ScanConf.scala 32:20]
  reg  confReg_516; // @[ScanConf.scala 32:20]
  reg  confReg_517; // @[ScanConf.scala 32:20]
  reg  confReg_518; // @[ScanConf.scala 32:20]
  reg  confReg_519; // @[ScanConf.scala 32:20]
  reg  confReg_520; // @[ScanConf.scala 32:20]
  reg  confReg_521; // @[ScanConf.scala 32:20]
  reg  confReg_522; // @[ScanConf.scala 32:20]
  reg  confReg_523; // @[ScanConf.scala 32:20]
  reg  confReg_524; // @[ScanConf.scala 32:20]
  reg  confReg_525; // @[ScanConf.scala 32:20]
  reg  confReg_526; // @[ScanConf.scala 32:20]
  reg  confReg_527; // @[ScanConf.scala 32:20]
  reg  confReg_528; // @[ScanConf.scala 32:20]
  reg  confReg_529; // @[ScanConf.scala 32:20]
  reg  confReg_530; // @[ScanConf.scala 32:20]
  reg  confReg_531; // @[ScanConf.scala 32:20]
  reg  confReg_532; // @[ScanConf.scala 32:20]
  reg  confReg_533; // @[ScanConf.scala 32:20]
  reg  confReg_534; // @[ScanConf.scala 32:20]
  reg  confReg_535; // @[ScanConf.scala 32:20]
  reg  confReg_536; // @[ScanConf.scala 32:20]
  reg  confReg_537; // @[ScanConf.scala 32:20]
  reg  confReg_538; // @[ScanConf.scala 32:20]
  reg  confReg_539; // @[ScanConf.scala 32:20]
  reg  confReg_540; // @[ScanConf.scala 32:20]
  reg  confReg_541; // @[ScanConf.scala 32:20]
  reg  confReg_542; // @[ScanConf.scala 32:20]
  reg  confReg_543; // @[ScanConf.scala 32:20]
  reg  confReg_544; // @[ScanConf.scala 32:20]
  reg  confReg_545; // @[ScanConf.scala 32:20]
  reg  confReg_546; // @[ScanConf.scala 32:20]
  reg  confReg_547; // @[ScanConf.scala 32:20]
  reg  confReg_548; // @[ScanConf.scala 32:20]
  reg  confReg_549; // @[ScanConf.scala 32:20]
  reg  confReg_550; // @[ScanConf.scala 32:20]
  reg  confReg_551; // @[ScanConf.scala 32:20]
  reg  confReg_552; // @[ScanConf.scala 32:20]
  reg  confReg_553; // @[ScanConf.scala 32:20]
  reg  confReg_554; // @[ScanConf.scala 32:20]
  reg  confReg_555; // @[ScanConf.scala 32:20]
  reg  confReg_556; // @[ScanConf.scala 32:20]
  reg  confReg_557; // @[ScanConf.scala 32:20]
  reg  confReg_558; // @[ScanConf.scala 32:20]
  reg  confReg_559; // @[ScanConf.scala 32:20]
  reg  confReg_560; // @[ScanConf.scala 32:20]
  reg  confReg_561; // @[ScanConf.scala 32:20]
  reg  confReg_562; // @[ScanConf.scala 32:20]
  reg  confReg_563; // @[ScanConf.scala 32:20]
  reg  confReg_564; // @[ScanConf.scala 32:20]
  reg  confReg_565; // @[ScanConf.scala 32:20]
  reg  confReg_566; // @[ScanConf.scala 32:20]
  reg  confReg_567; // @[ScanConf.scala 32:20]
  reg  confReg_568; // @[ScanConf.scala 32:20]
  reg  confReg_569; // @[ScanConf.scala 32:20]
  reg  confReg_570; // @[ScanConf.scala 32:20]
  reg  confReg_571; // @[ScanConf.scala 32:20]
  reg  confReg_572; // @[ScanConf.scala 32:20]
  reg  confReg_573; // @[ScanConf.scala 32:20]
  reg  confReg_574; // @[ScanConf.scala 32:20]
  reg  confReg_575; // @[ScanConf.scala 32:20]
  reg  confReg_576; // @[ScanConf.scala 32:20]
  reg  confReg_577; // @[ScanConf.scala 32:20]
  reg  confReg_578; // @[ScanConf.scala 32:20]
  reg  confReg_579; // @[ScanConf.scala 32:20]
  reg  confReg_580; // @[ScanConf.scala 32:20]
  reg  confReg_581; // @[ScanConf.scala 32:20]
  reg  confReg_582; // @[ScanConf.scala 32:20]
  reg  confReg_583; // @[ScanConf.scala 32:20]
  reg  confReg_584; // @[ScanConf.scala 32:20]
  reg  confReg_585; // @[ScanConf.scala 32:20]
  reg  confReg_586; // @[ScanConf.scala 32:20]
  reg  confReg_587; // @[ScanConf.scala 32:20]
  reg  confReg_588; // @[ScanConf.scala 32:20]
  reg  confReg_589; // @[ScanConf.scala 32:20]
  reg  confReg_590; // @[ScanConf.scala 32:20]
  reg  confReg_591; // @[ScanConf.scala 32:20]
  reg  confReg_592; // @[ScanConf.scala 32:20]
  reg  confReg_593; // @[ScanConf.scala 32:20]
  reg  confReg_594; // @[ScanConf.scala 32:20]
  reg  confReg_595; // @[ScanConf.scala 32:20]
  reg  confReg_596; // @[ScanConf.scala 32:20]
  reg  confReg_597; // @[ScanConf.scala 32:20]
  reg  confReg_598; // @[ScanConf.scala 32:20]
  reg  confReg_599; // @[ScanConf.scala 32:20]
  reg  confReg_600; // @[ScanConf.scala 32:20]
  reg  confReg_601; // @[ScanConf.scala 32:20]
  reg  confReg_602; // @[ScanConf.scala 32:20]
  reg  confReg_603; // @[ScanConf.scala 32:20]
  reg  confReg_604; // @[ScanConf.scala 32:20]
  reg  confReg_605; // @[ScanConf.scala 32:20]
  reg  confReg_606; // @[ScanConf.scala 32:20]
  reg  confReg_607; // @[ScanConf.scala 32:20]
  reg  confReg_608; // @[ScanConf.scala 32:20]
  reg  confReg_609; // @[ScanConf.scala 32:20]
  reg  confReg_610; // @[ScanConf.scala 32:20]
  reg  confReg_611; // @[ScanConf.scala 32:20]
  reg  confReg_612; // @[ScanConf.scala 32:20]
  reg  confReg_613; // @[ScanConf.scala 32:20]
  reg  confReg_614; // @[ScanConf.scala 32:20]
  reg  confReg_615; // @[ScanConf.scala 32:20]
  reg  confReg_616; // @[ScanConf.scala 32:20]
  reg  confReg_617; // @[ScanConf.scala 32:20]
  reg  confReg_618; // @[ScanConf.scala 32:20]
  reg  confReg_619; // @[ScanConf.scala 32:20]
  reg  confReg_620; // @[ScanConf.scala 32:20]
  reg  confReg_621; // @[ScanConf.scala 32:20]
  reg  confReg_622; // @[ScanConf.scala 32:20]
  reg  confReg_623; // @[ScanConf.scala 32:20]
  reg  confReg_624; // @[ScanConf.scala 32:20]
  reg  confReg_625; // @[ScanConf.scala 32:20]
  reg  confReg_626; // @[ScanConf.scala 32:20]
  reg  confReg_627; // @[ScanConf.scala 32:20]
  reg  confReg_628; // @[ScanConf.scala 32:20]
  reg  confReg_629; // @[ScanConf.scala 32:20]
  reg  confReg_630; // @[ScanConf.scala 32:20]
  reg  confReg_631; // @[ScanConf.scala 32:20]
  reg  confReg_632; // @[ScanConf.scala 32:20]
  reg  confReg_633; // @[ScanConf.scala 32:20]
  reg  confReg_634; // @[ScanConf.scala 32:20]
  reg  confReg_635; // @[ScanConf.scala 32:20]
  reg  confReg_636; // @[ScanConf.scala 32:20]
  reg  confReg_637; // @[ScanConf.scala 32:20]
  reg  confReg_638; // @[ScanConf.scala 32:20]
  reg  confReg_639; // @[ScanConf.scala 32:20]
  reg  confReg_640; // @[ScanConf.scala 32:20]
  reg  confReg_641; // @[ScanConf.scala 32:20]
  reg  confReg_642; // @[ScanConf.scala 32:20]
  reg  confReg_643; // @[ScanConf.scala 32:20]
  reg  confReg_644; // @[ScanConf.scala 32:20]
  reg  confReg_645; // @[ScanConf.scala 32:20]
  reg  confReg_646; // @[ScanConf.scala 32:20]
  reg  confReg_647; // @[ScanConf.scala 32:20]
  reg  confReg_648; // @[ScanConf.scala 32:20]
  reg  confReg_649; // @[ScanConf.scala 32:20]
  reg  confReg_650; // @[ScanConf.scala 32:20]
  reg  confReg_651; // @[ScanConf.scala 32:20]
  reg  confReg_652; // @[ScanConf.scala 32:20]
  reg  confReg_653; // @[ScanConf.scala 32:20]
  reg  confReg_654; // @[ScanConf.scala 32:20]
  reg  confReg_655; // @[ScanConf.scala 32:20]
  wire [7:0] io_scan_out_lo = {confReg_7,confReg_6,confReg_5,confReg_4,confReg_3,confReg_2,confReg_1,confReg_0}; // @[ScanConf.scala 46:47]
  wire [7:0] io_scan_out_hi = {confReg_15,confReg_14,confReg_13,confReg_12,confReg_11,confReg_10,confReg_9,confReg_8}; // @[ScanConf.scala 46:47]
  wire [9:0] io_confOut_lo_lo_lo_lo_lo_lo = {confReg_9,confReg_8,confReg_7,confReg_6,confReg_5,confReg_4,confReg_3,
    confReg_2,confReg_1,confReg_0}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_lo_lo_lo_hi = {confReg_19,confReg_18,confReg_17,confReg_16,confReg_15,confReg_14,
    confReg_13,confReg_12,confReg_11,confReg_10}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_lo_lo_hi_lo = {confReg_29,confReg_28,confReg_27,confReg_26,confReg_25,confReg_24,
    confReg_23,confReg_22,confReg_21,confReg_20}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_lo_lo_lo_lo_hi_hi_lo = {confReg_34,confReg_33,confReg_32,confReg_31,confReg_30}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_lo_lo_lo_lo = {confReg_40,confReg_39,confReg_38,confReg_37,confReg_36,confReg_35,
    io_confOut_lo_lo_lo_lo_hi_hi_lo,io_confOut_lo_lo_lo_lo_hi_lo,io_confOut_lo_lo_lo_lo_lo_hi,
    io_confOut_lo_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_lo_hi_lo_lo = {confReg_50,confReg_49,confReg_48,confReg_47,confReg_46,confReg_45,
    confReg_44,confReg_43,confReg_42,confReg_41}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_lo_hi_lo_hi = {confReg_60,confReg_59,confReg_58,confReg_57,confReg_56,confReg_55,
    confReg_54,confReg_53,confReg_52,confReg_51}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_lo_hi_hi_lo = {confReg_70,confReg_69,confReg_68,confReg_67,confReg_66,confReg_65,
    confReg_64,confReg_63,confReg_62,confReg_61}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_lo_lo_lo_hi_hi_hi_lo = {confReg_75,confReg_74,confReg_73,confReg_72,confReg_71}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_lo_lo_lo_hi = {confReg_81,confReg_80,confReg_79,confReg_78,confReg_77,confReg_76,
    io_confOut_lo_lo_lo_hi_hi_hi_lo,io_confOut_lo_lo_lo_hi_hi_lo,io_confOut_lo_lo_lo_hi_lo_hi,
    io_confOut_lo_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_hi_lo_lo_lo = {confReg_91,confReg_90,confReg_89,confReg_88,confReg_87,confReg_86,
    confReg_85,confReg_84,confReg_83,confReg_82}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_hi_lo_lo_hi = {confReg_101,confReg_100,confReg_99,confReg_98,confReg_97,confReg_96,
    confReg_95,confReg_94,confReg_93,confReg_92}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_hi_lo_hi_lo = {confReg_111,confReg_110,confReg_109,confReg_108,confReg_107,confReg_106,
    confReg_105,confReg_104,confReg_103,confReg_102}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_lo_lo_hi_lo_hi_hi_lo = {confReg_116,confReg_115,confReg_114,confReg_113,confReg_112}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_lo_lo_hi_lo = {confReg_122,confReg_121,confReg_120,confReg_119,confReg_118,confReg_117,
    io_confOut_lo_lo_hi_lo_hi_hi_lo,io_confOut_lo_lo_hi_lo_hi_lo,io_confOut_lo_lo_hi_lo_lo_hi,
    io_confOut_lo_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_hi_hi_lo_lo = {confReg_132,confReg_131,confReg_130,confReg_129,confReg_128,confReg_127,
    confReg_126,confReg_125,confReg_124,confReg_123}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_hi_hi_lo_hi = {confReg_142,confReg_141,confReg_140,confReg_139,confReg_138,confReg_137,
    confReg_136,confReg_135,confReg_134,confReg_133}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_lo_hi_hi_hi_lo = {confReg_152,confReg_151,confReg_150,confReg_149,confReg_148,confReg_147,
    confReg_146,confReg_145,confReg_144,confReg_143}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_lo_lo_hi_hi_hi_hi_lo = {confReg_157,confReg_156,confReg_155,confReg_154,confReg_153}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_lo_lo_hi_hi = {confReg_163,confReg_162,confReg_161,confReg_160,confReg_159,confReg_158,
    io_confOut_lo_lo_hi_hi_hi_hi_lo,io_confOut_lo_lo_hi_hi_hi_lo,io_confOut_lo_lo_hi_hi_lo_hi,
    io_confOut_lo_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_lo_lo_lo_lo = {confReg_173,confReg_172,confReg_171,confReg_170,confReg_169,confReg_168,
    confReg_167,confReg_166,confReg_165,confReg_164}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_lo_lo_lo_hi = {confReg_183,confReg_182,confReg_181,confReg_180,confReg_179,confReg_178,
    confReg_177,confReg_176,confReg_175,confReg_174}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_lo_lo_hi_lo = {confReg_193,confReg_192,confReg_191,confReg_190,confReg_189,confReg_188,
    confReg_187,confReg_186,confReg_185,confReg_184}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_lo_hi_lo_lo_hi_hi_lo = {confReg_198,confReg_197,confReg_196,confReg_195,confReg_194}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_lo_hi_lo_lo = {confReg_204,confReg_203,confReg_202,confReg_201,confReg_200,confReg_199,
    io_confOut_lo_hi_lo_lo_hi_hi_lo,io_confOut_lo_hi_lo_lo_hi_lo,io_confOut_lo_hi_lo_lo_lo_hi,
    io_confOut_lo_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_lo_hi_lo_lo = {confReg_214,confReg_213,confReg_212,confReg_211,confReg_210,confReg_209,
    confReg_208,confReg_207,confReg_206,confReg_205}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_lo_hi_lo_hi = {confReg_224,confReg_223,confReg_222,confReg_221,confReg_220,confReg_219,
    confReg_218,confReg_217,confReg_216,confReg_215}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_lo_hi_hi_lo = {confReg_234,confReg_233,confReg_232,confReg_231,confReg_230,confReg_229,
    confReg_228,confReg_227,confReg_226,confReg_225}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_lo_hi_lo_hi_hi_hi_lo = {confReg_239,confReg_238,confReg_237,confReg_236,confReg_235}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_lo_hi_lo_hi = {confReg_245,confReg_244,confReg_243,confReg_242,confReg_241,confReg_240,
    io_confOut_lo_hi_lo_hi_hi_hi_lo,io_confOut_lo_hi_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi_lo_hi,
    io_confOut_lo_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_hi_lo_lo_lo = {confReg_255,confReg_254,confReg_253,confReg_252,confReg_251,confReg_250,
    confReg_249,confReg_248,confReg_247,confReg_246}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_hi_lo_lo_hi = {confReg_265,confReg_264,confReg_263,confReg_262,confReg_261,confReg_260,
    confReg_259,confReg_258,confReg_257,confReg_256}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_hi_lo_hi_lo = {confReg_275,confReg_274,confReg_273,confReg_272,confReg_271,confReg_270,
    confReg_269,confReg_268,confReg_267,confReg_266}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_lo_hi_hi_lo_hi_hi_lo = {confReg_280,confReg_279,confReg_278,confReg_277,confReg_276}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_lo_hi_hi_lo = {confReg_286,confReg_285,confReg_284,confReg_283,confReg_282,confReg_281,
    io_confOut_lo_hi_hi_lo_hi_hi_lo,io_confOut_lo_hi_hi_lo_hi_lo,io_confOut_lo_hi_hi_lo_lo_hi,
    io_confOut_lo_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_hi_hi_lo_lo = {confReg_296,confReg_295,confReg_294,confReg_293,confReg_292,confReg_291,
    confReg_290,confReg_289,confReg_288,confReg_287}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_hi_hi_lo_hi = {confReg_306,confReg_305,confReg_304,confReg_303,confReg_302,confReg_301,
    confReg_300,confReg_299,confReg_298,confReg_297}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_lo_hi_hi_hi_hi_lo = {confReg_316,confReg_315,confReg_314,confReg_313,confReg_312,confReg_311,
    confReg_310,confReg_309,confReg_308,confReg_307}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_lo_hi_hi_hi_hi_hi_lo = {confReg_321,confReg_320,confReg_319,confReg_318,confReg_317}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_lo_hi_hi_hi = {confReg_327,confReg_326,confReg_325,confReg_324,confReg_323,confReg_322,
    io_confOut_lo_hi_hi_hi_hi_hi_lo,io_confOut_lo_hi_hi_hi_hi_lo,io_confOut_lo_hi_hi_hi_lo_hi,
    io_confOut_lo_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [327:0] io_confOut_lo = {io_confOut_lo_hi_hi_hi,io_confOut_lo_hi_hi_lo,io_confOut_lo_hi_lo_hi,
    io_confOut_lo_hi_lo_lo,io_confOut_lo_lo_hi_hi,io_confOut_lo_lo_hi_lo,io_confOut_lo_lo_lo_hi,io_confOut_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_lo_lo_lo_lo = {confReg_337,confReg_336,confReg_335,confReg_334,confReg_333,confReg_332,
    confReg_331,confReg_330,confReg_329,confReg_328}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_lo_lo_lo_hi = {confReg_347,confReg_346,confReg_345,confReg_344,confReg_343,confReg_342,
    confReg_341,confReg_340,confReg_339,confReg_338}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_lo_lo_hi_lo = {confReg_357,confReg_356,confReg_355,confReg_354,confReg_353,confReg_352,
    confReg_351,confReg_350,confReg_349,confReg_348}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_hi_lo_lo_lo_hi_hi_lo = {confReg_362,confReg_361,confReg_360,confReg_359,confReg_358}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_hi_lo_lo_lo = {confReg_368,confReg_367,confReg_366,confReg_365,confReg_364,confReg_363,
    io_confOut_hi_lo_lo_lo_hi_hi_lo,io_confOut_hi_lo_lo_lo_hi_lo,io_confOut_hi_lo_lo_lo_lo_hi,
    io_confOut_hi_lo_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_lo_hi_lo_lo = {confReg_378,confReg_377,confReg_376,confReg_375,confReg_374,confReg_373,
    confReg_372,confReg_371,confReg_370,confReg_369}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_lo_hi_lo_hi = {confReg_388,confReg_387,confReg_386,confReg_385,confReg_384,confReg_383,
    confReg_382,confReg_381,confReg_380,confReg_379}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_lo_hi_hi_lo = {confReg_398,confReg_397,confReg_396,confReg_395,confReg_394,confReg_393,
    confReg_392,confReg_391,confReg_390,confReg_389}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_hi_lo_lo_hi_hi_hi_lo = {confReg_403,confReg_402,confReg_401,confReg_400,confReg_399}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_hi_lo_lo_hi = {confReg_409,confReg_408,confReg_407,confReg_406,confReg_405,confReg_404,
    io_confOut_hi_lo_lo_hi_hi_hi_lo,io_confOut_hi_lo_lo_hi_hi_lo,io_confOut_hi_lo_lo_hi_lo_hi,
    io_confOut_hi_lo_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_hi_lo_lo_lo = {confReg_419,confReg_418,confReg_417,confReg_416,confReg_415,confReg_414,
    confReg_413,confReg_412,confReg_411,confReg_410}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_hi_lo_lo_hi = {confReg_429,confReg_428,confReg_427,confReg_426,confReg_425,confReg_424,
    confReg_423,confReg_422,confReg_421,confReg_420}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_hi_lo_hi_lo = {confReg_439,confReg_438,confReg_437,confReg_436,confReg_435,confReg_434,
    confReg_433,confReg_432,confReg_431,confReg_430}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_hi_lo_hi_lo_hi_hi_lo = {confReg_444,confReg_443,confReg_442,confReg_441,confReg_440}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_hi_lo_hi_lo = {confReg_450,confReg_449,confReg_448,confReg_447,confReg_446,confReg_445,
    io_confOut_hi_lo_hi_lo_hi_hi_lo,io_confOut_hi_lo_hi_lo_hi_lo,io_confOut_hi_lo_hi_lo_lo_hi,
    io_confOut_hi_lo_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_hi_hi_lo_lo = {confReg_460,confReg_459,confReg_458,confReg_457,confReg_456,confReg_455,
    confReg_454,confReg_453,confReg_452,confReg_451}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_hi_hi_lo_hi = {confReg_470,confReg_469,confReg_468,confReg_467,confReg_466,confReg_465,
    confReg_464,confReg_463,confReg_462,confReg_461}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_lo_hi_hi_hi_lo = {confReg_480,confReg_479,confReg_478,confReg_477,confReg_476,confReg_475,
    confReg_474,confReg_473,confReg_472,confReg_471}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_hi_lo_hi_hi_hi_hi_lo = {confReg_485,confReg_484,confReg_483,confReg_482,confReg_481}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_hi_lo_hi_hi = {confReg_491,confReg_490,confReg_489,confReg_488,confReg_487,confReg_486,
    io_confOut_hi_lo_hi_hi_hi_hi_lo,io_confOut_hi_lo_hi_hi_hi_lo,io_confOut_hi_lo_hi_hi_lo_hi,
    io_confOut_hi_lo_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_lo_lo_lo_lo = {confReg_501,confReg_500,confReg_499,confReg_498,confReg_497,confReg_496,
    confReg_495,confReg_494,confReg_493,confReg_492}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_lo_lo_lo_hi = {confReg_511,confReg_510,confReg_509,confReg_508,confReg_507,confReg_506,
    confReg_505,confReg_504,confReg_503,confReg_502}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_lo_lo_hi_lo = {confReg_521,confReg_520,confReg_519,confReg_518,confReg_517,confReg_516,
    confReg_515,confReg_514,confReg_513,confReg_512}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_hi_hi_lo_lo_hi_hi_lo = {confReg_526,confReg_525,confReg_524,confReg_523,confReg_522}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_hi_hi_lo_lo = {confReg_532,confReg_531,confReg_530,confReg_529,confReg_528,confReg_527,
    io_confOut_hi_hi_lo_lo_hi_hi_lo,io_confOut_hi_hi_lo_lo_hi_lo,io_confOut_hi_hi_lo_lo_lo_hi,
    io_confOut_hi_hi_lo_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_lo_hi_lo_lo = {confReg_542,confReg_541,confReg_540,confReg_539,confReg_538,confReg_537,
    confReg_536,confReg_535,confReg_534,confReg_533}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_lo_hi_lo_hi = {confReg_552,confReg_551,confReg_550,confReg_549,confReg_548,confReg_547,
    confReg_546,confReg_545,confReg_544,confReg_543}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_lo_hi_hi_lo = {confReg_562,confReg_561,confReg_560,confReg_559,confReg_558,confReg_557,
    confReg_556,confReg_555,confReg_554,confReg_553}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_hi_hi_lo_hi_hi_hi_lo = {confReg_567,confReg_566,confReg_565,confReg_564,confReg_563}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_hi_hi_lo_hi = {confReg_573,confReg_572,confReg_571,confReg_570,confReg_569,confReg_568,
    io_confOut_hi_hi_lo_hi_hi_hi_lo,io_confOut_hi_hi_lo_hi_hi_lo,io_confOut_hi_hi_lo_hi_lo_hi,
    io_confOut_hi_hi_lo_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_hi_lo_lo_lo = {confReg_583,confReg_582,confReg_581,confReg_580,confReg_579,confReg_578,
    confReg_577,confReg_576,confReg_575,confReg_574}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_hi_lo_lo_hi = {confReg_593,confReg_592,confReg_591,confReg_590,confReg_589,confReg_588,
    confReg_587,confReg_586,confReg_585,confReg_584}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_hi_lo_hi_lo = {confReg_603,confReg_602,confReg_601,confReg_600,confReg_599,confReg_598,
    confReg_597,confReg_596,confReg_595,confReg_594}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_hi_hi_hi_lo_hi_hi_lo = {confReg_608,confReg_607,confReg_606,confReg_605,confReg_604}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_hi_hi_hi_lo = {confReg_614,confReg_613,confReg_612,confReg_611,confReg_610,confReg_609,
    io_confOut_hi_hi_hi_lo_hi_hi_lo,io_confOut_hi_hi_hi_lo_hi_lo,io_confOut_hi_hi_hi_lo_lo_hi,
    io_confOut_hi_hi_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_hi_hi_lo_lo = {confReg_624,confReg_623,confReg_622,confReg_621,confReg_620,confReg_619,
    confReg_618,confReg_617,confReg_616,confReg_615}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_hi_hi_lo_hi = {confReg_634,confReg_633,confReg_632,confReg_631,confReg_630,confReg_629,
    confReg_628,confReg_627,confReg_626,confReg_625}; // @[ScanConf.scala 48:25]
  wire [9:0] io_confOut_hi_hi_hi_hi_hi_lo = {confReg_644,confReg_643,confReg_642,confReg_641,confReg_640,confReg_639,
    confReg_638,confReg_637,confReg_636,confReg_635}; // @[ScanConf.scala 48:25]
  wire [4:0] io_confOut_hi_hi_hi_hi_hi_hi_lo = {confReg_649,confReg_648,confReg_647,confReg_646,confReg_645}; // @[ScanConf.scala 48:25]
  wire [40:0] io_confOut_hi_hi_hi_hi = {confReg_655,confReg_654,confReg_653,confReg_652,confReg_651,confReg_650,
    io_confOut_hi_hi_hi_hi_hi_hi_lo,io_confOut_hi_hi_hi_hi_hi_lo,io_confOut_hi_hi_hi_hi_lo_hi,
    io_confOut_hi_hi_hi_hi_lo_lo}; // @[ScanConf.scala 48:25]
  wire [327:0] io_confOut_hi = {io_confOut_hi_hi_hi_hi,io_confOut_hi_hi_hi_lo,io_confOut_hi_hi_lo_hi,
    io_confOut_hi_hi_lo_lo,io_confOut_hi_lo_hi_hi,io_confOut_hi_lo_hi_lo,io_confOut_hi_lo_lo_hi,io_confOut_hi_lo_lo_lo}; // @[ScanConf.scala 48:25]
  assign ioBundle_confOut = {io_confOut_hi,io_confOut_lo}; // @[ScanConf.scala 48:25]
  assign ioBundle_scan_out = {io_scan_out_hi,io_scan_out_lo}; // @[ScanConf.scala 46:47]
  always @(posedge clock) begin
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_0 <= confReg_16; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_1 <= confReg_17; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_2 <= confReg_18; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_3 <= confReg_19; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_4 <= confReg_20; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_5 <= confReg_21; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_6 <= confReg_22; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_7 <= confReg_23; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_8 <= confReg_24; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_9 <= confReg_25; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_10 <= confReg_26; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_11 <= confReg_27; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_12 <= confReg_28; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_13 <= confReg_29; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_14 <= confReg_30; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_15 <= confReg_31; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_16 <= confReg_32; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_17 <= confReg_33; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_18 <= confReg_34; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_19 <= confReg_35; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_20 <= confReg_36; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_21 <= confReg_37; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_22 <= confReg_38; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_23 <= confReg_39; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_24 <= confReg_40; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_25 <= confReg_41; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_26 <= confReg_42; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_27 <= confReg_43; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_28 <= confReg_44; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_29 <= confReg_45; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_30 <= confReg_46; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_31 <= confReg_47; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_32 <= confReg_48; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_33 <= confReg_49; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_34 <= confReg_50; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_35 <= confReg_51; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_36 <= confReg_52; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_37 <= confReg_53; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_38 <= confReg_54; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_39 <= confReg_55; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_40 <= confReg_56; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_41 <= confReg_57; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_42 <= confReg_58; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_43 <= confReg_59; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_44 <= confReg_60; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_45 <= confReg_61; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_46 <= confReg_62; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_47 <= confReg_63; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_48 <= confReg_64; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_49 <= confReg_65; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_50 <= confReg_66; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_51 <= confReg_67; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_52 <= confReg_68; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_53 <= confReg_69; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_54 <= confReg_70; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_55 <= confReg_71; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_56 <= confReg_72; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_57 <= confReg_73; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_58 <= confReg_74; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_59 <= confReg_75; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_60 <= confReg_76; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_61 <= confReg_77; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_62 <= confReg_78; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_63 <= confReg_79; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_64 <= confReg_80; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_65 <= confReg_81; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_66 <= confReg_82; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_67 <= confReg_83; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_68 <= confReg_84; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_69 <= confReg_85; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_70 <= confReg_86; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_71 <= confReg_87; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_72 <= confReg_88; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_73 <= confReg_89; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_74 <= confReg_90; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_75 <= confReg_91; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_76 <= confReg_92; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_77 <= confReg_93; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_78 <= confReg_94; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_79 <= confReg_95; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_80 <= confReg_96; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_81 <= confReg_97; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_82 <= confReg_98; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_83 <= confReg_99; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_84 <= confReg_100; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_85 <= confReg_101; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_86 <= confReg_102; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_87 <= confReg_103; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_88 <= confReg_104; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_89 <= confReg_105; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_90 <= confReg_106; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_91 <= confReg_107; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_92 <= confReg_108; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_93 <= confReg_109; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_94 <= confReg_110; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_95 <= confReg_111; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_96 <= confReg_112; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_97 <= confReg_113; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_98 <= confReg_114; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_99 <= confReg_115; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_100 <= confReg_116; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_101 <= confReg_117; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_102 <= confReg_118; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_103 <= confReg_119; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_104 <= confReg_120; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_105 <= confReg_121; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_106 <= confReg_122; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_107 <= confReg_123; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_108 <= confReg_124; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_109 <= confReg_125; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_110 <= confReg_126; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_111 <= confReg_127; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_112 <= confReg_128; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_113 <= confReg_129; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_114 <= confReg_130; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_115 <= confReg_131; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_116 <= confReg_132; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_117 <= confReg_133; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_118 <= confReg_134; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_119 <= confReg_135; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_120 <= confReg_136; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_121 <= confReg_137; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_122 <= confReg_138; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_123 <= confReg_139; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_124 <= confReg_140; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_125 <= confReg_141; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_126 <= confReg_142; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_127 <= confReg_143; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_128 <= confReg_144; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_129 <= confReg_145; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_130 <= confReg_146; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_131 <= confReg_147; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_132 <= confReg_148; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_133 <= confReg_149; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_134 <= confReg_150; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_135 <= confReg_151; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_136 <= confReg_152; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_137 <= confReg_153; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_138 <= confReg_154; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_139 <= confReg_155; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_140 <= confReg_156; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_141 <= confReg_157; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_142 <= confReg_158; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_143 <= confReg_159; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_144 <= confReg_160; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_145 <= confReg_161; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_146 <= confReg_162; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_147 <= confReg_163; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_148 <= confReg_164; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_149 <= confReg_165; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_150 <= confReg_166; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_151 <= confReg_167; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_152 <= confReg_168; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_153 <= confReg_169; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_154 <= confReg_170; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_155 <= confReg_171; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_156 <= confReg_172; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_157 <= confReg_173; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_158 <= confReg_174; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_159 <= confReg_175; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_160 <= confReg_176; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_161 <= confReg_177; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_162 <= confReg_178; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_163 <= confReg_179; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_164 <= confReg_180; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_165 <= confReg_181; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_166 <= confReg_182; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_167 <= confReg_183; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_168 <= confReg_184; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_169 <= confReg_185; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_170 <= confReg_186; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_171 <= confReg_187; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_172 <= confReg_188; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_173 <= confReg_189; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_174 <= confReg_190; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_175 <= confReg_191; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_176 <= confReg_192; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_177 <= confReg_193; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_178 <= confReg_194; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_179 <= confReg_195; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_180 <= confReg_196; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_181 <= confReg_197; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_182 <= confReg_198; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_183 <= confReg_199; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_184 <= confReg_200; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_185 <= confReg_201; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_186 <= confReg_202; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_187 <= confReg_203; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_188 <= confReg_204; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_189 <= confReg_205; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_190 <= confReg_206; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_191 <= confReg_207; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_192 <= confReg_208; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_193 <= confReg_209; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_194 <= confReg_210; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_195 <= confReg_211; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_196 <= confReg_212; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_197 <= confReg_213; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_198 <= confReg_214; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_199 <= confReg_215; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_200 <= confReg_216; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_201 <= confReg_217; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_202 <= confReg_218; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_203 <= confReg_219; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_204 <= confReg_220; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_205 <= confReg_221; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_206 <= confReg_222; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_207 <= confReg_223; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_208 <= confReg_224; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_209 <= confReg_225; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_210 <= confReg_226; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_211 <= confReg_227; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_212 <= confReg_228; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_213 <= confReg_229; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_214 <= confReg_230; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_215 <= confReg_231; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_216 <= confReg_232; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_217 <= confReg_233; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_218 <= confReg_234; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_219 <= confReg_235; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_220 <= confReg_236; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_221 <= confReg_237; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_222 <= confReg_238; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_223 <= confReg_239; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_224 <= confReg_240; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_225 <= confReg_241; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_226 <= confReg_242; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_227 <= confReg_243; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_228 <= confReg_244; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_229 <= confReg_245; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_230 <= confReg_246; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_231 <= confReg_247; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_232 <= confReg_248; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_233 <= confReg_249; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_234 <= confReg_250; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_235 <= confReg_251; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_236 <= confReg_252; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_237 <= confReg_253; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_238 <= confReg_254; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_239 <= confReg_255; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_240 <= confReg_256; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_241 <= confReg_257; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_242 <= confReg_258; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_243 <= confReg_259; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_244 <= confReg_260; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_245 <= confReg_261; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_246 <= confReg_262; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_247 <= confReg_263; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_248 <= confReg_264; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_249 <= confReg_265; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_250 <= confReg_266; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_251 <= confReg_267; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_252 <= confReg_268; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_253 <= confReg_269; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_254 <= confReg_270; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_255 <= confReg_271; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_256 <= confReg_272; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_257 <= confReg_273; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_258 <= confReg_274; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_259 <= confReg_275; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_260 <= confReg_276; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_261 <= confReg_277; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_262 <= confReg_278; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_263 <= confReg_279; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_264 <= confReg_280; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_265 <= confReg_281; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_266 <= confReg_282; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_267 <= confReg_283; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_268 <= confReg_284; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_269 <= confReg_285; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_270 <= confReg_286; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_271 <= confReg_287; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_272 <= confReg_288; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_273 <= confReg_289; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_274 <= confReg_290; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_275 <= confReg_291; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_276 <= confReg_292; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_277 <= confReg_293; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_278 <= confReg_294; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_279 <= confReg_295; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_280 <= confReg_296; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_281 <= confReg_297; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_282 <= confReg_298; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_283 <= confReg_299; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_284 <= confReg_300; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_285 <= confReg_301; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_286 <= confReg_302; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_287 <= confReg_303; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_288 <= confReg_304; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_289 <= confReg_305; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_290 <= confReg_306; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_291 <= confReg_307; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_292 <= confReg_308; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_293 <= confReg_309; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_294 <= confReg_310; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_295 <= confReg_311; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_296 <= confReg_312; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_297 <= confReg_313; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_298 <= confReg_314; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_299 <= confReg_315; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_300 <= confReg_316; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_301 <= confReg_317; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_302 <= confReg_318; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_303 <= confReg_319; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_304 <= confReg_320; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_305 <= confReg_321; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_306 <= confReg_322; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_307 <= confReg_323; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_308 <= confReg_324; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_309 <= confReg_325; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_310 <= confReg_326; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_311 <= confReg_327; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_312 <= confReg_328; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_313 <= confReg_329; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_314 <= confReg_330; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_315 <= confReg_331; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_316 <= confReg_332; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_317 <= confReg_333; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_318 <= confReg_334; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_319 <= confReg_335; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_320 <= confReg_336; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_321 <= confReg_337; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_322 <= confReg_338; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_323 <= confReg_339; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_324 <= confReg_340; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_325 <= confReg_341; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_326 <= confReg_342; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_327 <= confReg_343; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_328 <= confReg_344; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_329 <= confReg_345; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_330 <= confReg_346; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_331 <= confReg_347; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_332 <= confReg_348; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_333 <= confReg_349; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_334 <= confReg_350; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_335 <= confReg_351; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_336 <= confReg_352; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_337 <= confReg_353; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_338 <= confReg_354; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_339 <= confReg_355; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_340 <= confReg_356; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_341 <= confReg_357; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_342 <= confReg_358; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_343 <= confReg_359; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_344 <= confReg_360; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_345 <= confReg_361; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_346 <= confReg_362; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_347 <= confReg_363; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_348 <= confReg_364; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_349 <= confReg_365; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_350 <= confReg_366; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_351 <= confReg_367; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_352 <= confReg_368; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_353 <= confReg_369; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_354 <= confReg_370; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_355 <= confReg_371; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_356 <= confReg_372; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_357 <= confReg_373; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_358 <= confReg_374; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_359 <= confReg_375; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_360 <= confReg_376; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_361 <= confReg_377; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_362 <= confReg_378; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_363 <= confReg_379; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_364 <= confReg_380; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_365 <= confReg_381; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_366 <= confReg_382; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_367 <= confReg_383; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_368 <= confReg_384; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_369 <= confReg_385; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_370 <= confReg_386; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_371 <= confReg_387; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_372 <= confReg_388; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_373 <= confReg_389; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_374 <= confReg_390; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_375 <= confReg_391; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_376 <= confReg_392; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_377 <= confReg_393; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_378 <= confReg_394; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_379 <= confReg_395; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_380 <= confReg_396; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_381 <= confReg_397; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_382 <= confReg_398; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_383 <= confReg_399; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_384 <= confReg_400; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_385 <= confReg_401; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_386 <= confReg_402; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_387 <= confReg_403; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_388 <= confReg_404; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_389 <= confReg_405; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_390 <= confReg_406; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_391 <= confReg_407; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_392 <= confReg_408; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_393 <= confReg_409; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_394 <= confReg_410; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_395 <= confReg_411; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_396 <= confReg_412; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_397 <= confReg_413; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_398 <= confReg_414; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_399 <= confReg_415; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_400 <= confReg_416; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_401 <= confReg_417; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_402 <= confReg_418; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_403 <= confReg_419; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_404 <= confReg_420; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_405 <= confReg_421; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_406 <= confReg_422; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_407 <= confReg_423; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_408 <= confReg_424; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_409 <= confReg_425; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_410 <= confReg_426; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_411 <= confReg_427; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_412 <= confReg_428; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_413 <= confReg_429; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_414 <= confReg_430; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_415 <= confReg_431; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_416 <= confReg_432; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_417 <= confReg_433; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_418 <= confReg_434; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_419 <= confReg_435; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_420 <= confReg_436; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_421 <= confReg_437; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_422 <= confReg_438; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_423 <= confReg_439; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_424 <= confReg_440; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_425 <= confReg_441; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_426 <= confReg_442; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_427 <= confReg_443; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_428 <= confReg_444; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_429 <= confReg_445; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_430 <= confReg_446; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_431 <= confReg_447; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_432 <= confReg_448; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_433 <= confReg_449; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_434 <= confReg_450; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_435 <= confReg_451; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_436 <= confReg_452; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_437 <= confReg_453; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_438 <= confReg_454; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_439 <= confReg_455; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_440 <= confReg_456; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_441 <= confReg_457; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_442 <= confReg_458; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_443 <= confReg_459; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_444 <= confReg_460; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_445 <= confReg_461; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_446 <= confReg_462; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_447 <= confReg_463; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_448 <= confReg_464; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_449 <= confReg_465; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_450 <= confReg_466; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_451 <= confReg_467; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_452 <= confReg_468; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_453 <= confReg_469; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_454 <= confReg_470; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_455 <= confReg_471; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_456 <= confReg_472; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_457 <= confReg_473; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_458 <= confReg_474; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_459 <= confReg_475; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_460 <= confReg_476; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_461 <= confReg_477; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_462 <= confReg_478; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_463 <= confReg_479; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_464 <= confReg_480; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_465 <= confReg_481; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_466 <= confReg_482; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_467 <= confReg_483; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_468 <= confReg_484; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_469 <= confReg_485; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_470 <= confReg_486; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_471 <= confReg_487; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_472 <= confReg_488; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_473 <= confReg_489; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_474 <= confReg_490; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_475 <= confReg_491; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_476 <= confReg_492; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_477 <= confReg_493; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_478 <= confReg_494; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_479 <= confReg_495; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_480 <= confReg_496; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_481 <= confReg_497; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_482 <= confReg_498; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_483 <= confReg_499; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_484 <= confReg_500; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_485 <= confReg_501; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_486 <= confReg_502; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_487 <= confReg_503; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_488 <= confReg_504; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_489 <= confReg_505; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_490 <= confReg_506; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_491 <= confReg_507; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_492 <= confReg_508; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_493 <= confReg_509; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_494 <= confReg_510; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_495 <= confReg_511; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_496 <= confReg_512; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_497 <= confReg_513; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_498 <= confReg_514; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_499 <= confReg_515; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_500 <= confReg_516; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_501 <= confReg_517; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_502 <= confReg_518; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_503 <= confReg_519; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_504 <= confReg_520; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_505 <= confReg_521; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_506 <= confReg_522; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_507 <= confReg_523; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_508 <= confReg_524; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_509 <= confReg_525; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_510 <= confReg_526; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_511 <= confReg_527; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_512 <= confReg_528; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_513 <= confReg_529; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_514 <= confReg_530; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_515 <= confReg_531; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_516 <= confReg_532; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_517 <= confReg_533; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_518 <= confReg_534; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_519 <= confReg_535; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_520 <= confReg_536; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_521 <= confReg_537; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_522 <= confReg_538; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_523 <= confReg_539; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_524 <= confReg_540; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_525 <= confReg_541; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_526 <= confReg_542; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_527 <= confReg_543; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_528 <= confReg_544; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_529 <= confReg_545; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_530 <= confReg_546; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_531 <= confReg_547; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_532 <= confReg_548; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_533 <= confReg_549; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_534 <= confReg_550; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_535 <= confReg_551; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_536 <= confReg_552; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_537 <= confReg_553; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_538 <= confReg_554; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_539 <= confReg_555; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_540 <= confReg_556; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_541 <= confReg_557; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_542 <= confReg_558; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_543 <= confReg_559; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_544 <= confReg_560; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_545 <= confReg_561; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_546 <= confReg_562; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_547 <= confReg_563; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_548 <= confReg_564; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_549 <= confReg_565; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_550 <= confReg_566; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_551 <= confReg_567; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_552 <= confReg_568; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_553 <= confReg_569; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_554 <= confReg_570; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_555 <= confReg_571; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_556 <= confReg_572; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_557 <= confReg_573; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_558 <= confReg_574; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_559 <= confReg_575; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_560 <= confReg_576; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_561 <= confReg_577; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_562 <= confReg_578; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_563 <= confReg_579; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_564 <= confReg_580; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_565 <= confReg_581; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_566 <= confReg_582; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_567 <= confReg_583; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_568 <= confReg_584; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_569 <= confReg_585; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_570 <= confReg_586; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_571 <= confReg_587; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_572 <= confReg_588; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_573 <= confReg_589; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_574 <= confReg_590; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_575 <= confReg_591; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_576 <= confReg_592; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_577 <= confReg_593; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_578 <= confReg_594; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_579 <= confReg_595; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_580 <= confReg_596; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_581 <= confReg_597; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_582 <= confReg_598; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_583 <= confReg_599; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_584 <= confReg_600; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_585 <= confReg_601; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_586 <= confReg_602; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_587 <= confReg_603; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_588 <= confReg_604; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_589 <= confReg_605; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_590 <= confReg_606; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_591 <= confReg_607; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_592 <= confReg_608; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_593 <= confReg_609; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_594 <= confReg_610; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_595 <= confReg_611; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_596 <= confReg_612; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_597 <= confReg_613; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_598 <= confReg_614; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_599 <= confReg_615; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_600 <= confReg_616; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_601 <= confReg_617; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_602 <= confReg_618; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_603 <= confReg_619; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_604 <= confReg_620; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_605 <= confReg_621; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_606 <= confReg_622; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_607 <= confReg_623; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_608 <= confReg_624; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_609 <= confReg_625; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_610 <= confReg_626; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_611 <= confReg_627; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_612 <= confReg_628; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_613 <= confReg_629; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_614 <= confReg_630; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_615 <= confReg_631; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_616 <= confReg_632; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_617 <= confReg_633; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_618 <= confReg_634; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_619 <= confReg_635; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_620 <= confReg_636; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_621 <= confReg_637; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_622 <= confReg_638; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_623 <= confReg_639; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_624 <= confReg_640; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_625 <= confReg_641; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_626 <= confReg_642; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_627 <= confReg_643; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_628 <= confReg_644; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_629 <= confReg_645; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_630 <= confReg_646; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_631 <= confReg_647; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_632 <= confReg_648; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_633 <= confReg_649; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_634 <= confReg_650; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_635 <= confReg_651; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_636 <= confReg_652; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_637 <= confReg_653; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_638 <= confReg_654; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_639 <= confReg_655; // @[ScanConf.scala 41:36]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_640 <= ioBundle_scan_in[0]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_641 <= ioBundle_scan_in[1]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_642 <= ioBundle_scan_in[2]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_643 <= ioBundle_scan_in[3]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_644 <= ioBundle_scan_in[4]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_645 <= ioBundle_scan_in[5]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_646 <= ioBundle_scan_in[6]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_647 <= ioBundle_scan_in[7]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_648 <= ioBundle_scan_in[8]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_649 <= ioBundle_scan_in[9]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_650 <= ioBundle_scan_in[10]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_651 <= ioBundle_scan_in[11]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_652 <= ioBundle_scan_in[12]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_653 <= ioBundle_scan_in[13]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_654 <= ioBundle_scan_in[14]; // @[ScanConf.scala 38:72]
    end
    if (ioBundle_scan_en) begin // @[ScanConf.scala 37:20]
      confReg_655 <= ioBundle_scan_in[15]; // @[ScanConf.scala 38:72]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  confReg_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  confReg_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  confReg_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  confReg_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  confReg_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  confReg_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  confReg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  confReg_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  confReg_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  confReg_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  confReg_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  confReg_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  confReg_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  confReg_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  confReg_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  confReg_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  confReg_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  confReg_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  confReg_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  confReg_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  confReg_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  confReg_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  confReg_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  confReg_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  confReg_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  confReg_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  confReg_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  confReg_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  confReg_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  confReg_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  confReg_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  confReg_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  confReg_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  confReg_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  confReg_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  confReg_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  confReg_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  confReg_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  confReg_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  confReg_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  confReg_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  confReg_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  confReg_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  confReg_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  confReg_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  confReg_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  confReg_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  confReg_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  confReg_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  confReg_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  confReg_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  confReg_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  confReg_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  confReg_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  confReg_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  confReg_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  confReg_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  confReg_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  confReg_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  confReg_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  confReg_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  confReg_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  confReg_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  confReg_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  confReg_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  confReg_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  confReg_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  confReg_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  confReg_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  confReg_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  confReg_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  confReg_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  confReg_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  confReg_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  confReg_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  confReg_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  confReg_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  confReg_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  confReg_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  confReg_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  confReg_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  confReg_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  confReg_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  confReg_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  confReg_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  confReg_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  confReg_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  confReg_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  confReg_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  confReg_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  confReg_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  confReg_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  confReg_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  confReg_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  confReg_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  confReg_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  confReg_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  confReg_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  confReg_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  confReg_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  confReg_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  confReg_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  confReg_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  confReg_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  confReg_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  confReg_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  confReg_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  confReg_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  confReg_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  confReg_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  confReg_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  confReg_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  confReg_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  confReg_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  confReg_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  confReg_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  confReg_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  confReg_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  confReg_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  confReg_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  confReg_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  confReg_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  confReg_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  confReg_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  confReg_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  confReg_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  confReg_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  confReg_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  confReg_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  confReg_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  confReg_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  confReg_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  confReg_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  confReg_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  confReg_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  confReg_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  confReg_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  confReg_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  confReg_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  confReg_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  confReg_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  confReg_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  confReg_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  confReg_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  confReg_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  confReg_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  confReg_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  confReg_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  confReg_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  confReg_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  confReg_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  confReg_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  confReg_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  confReg_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  confReg_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  confReg_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  confReg_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  confReg_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  confReg_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  confReg_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  confReg_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  confReg_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  confReg_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  confReg_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  confReg_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  confReg_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  confReg_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  confReg_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  confReg_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  confReg_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  confReg_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  confReg_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  confReg_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  confReg_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  confReg_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  confReg_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  confReg_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  confReg_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  confReg_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  confReg_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  confReg_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  confReg_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  confReg_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  confReg_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  confReg_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  confReg_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  confReg_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  confReg_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  confReg_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  confReg_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  confReg_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  confReg_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  confReg_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  confReg_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  confReg_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  confReg_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  confReg_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  confReg_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  confReg_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  confReg_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  confReg_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  confReg_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  confReg_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  confReg_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  confReg_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  confReg_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  confReg_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  confReg_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  confReg_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  confReg_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  confReg_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  confReg_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  confReg_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  confReg_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  confReg_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  confReg_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  confReg_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  confReg_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  confReg_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  confReg_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  confReg_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  confReg_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  confReg_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  confReg_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  confReg_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  confReg_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  confReg_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  confReg_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  confReg_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  confReg_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  confReg_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  confReg_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  confReg_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  confReg_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  confReg_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  confReg_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  confReg_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  confReg_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  confReg_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  confReg_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  confReg_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  confReg_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  confReg_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  confReg_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  confReg_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  confReg_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  confReg_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  confReg_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  confReg_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  confReg_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  confReg_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  confReg_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  confReg_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  confReg_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  confReg_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  confReg_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  confReg_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  confReg_257 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  confReg_258 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  confReg_259 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  confReg_260 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  confReg_261 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  confReg_262 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  confReg_263 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  confReg_264 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  confReg_265 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  confReg_266 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  confReg_267 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  confReg_268 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  confReg_269 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  confReg_270 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  confReg_271 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  confReg_272 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  confReg_273 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  confReg_274 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  confReg_275 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  confReg_276 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  confReg_277 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  confReg_278 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  confReg_279 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  confReg_280 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  confReg_281 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  confReg_282 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  confReg_283 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  confReg_284 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  confReg_285 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  confReg_286 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  confReg_287 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  confReg_288 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  confReg_289 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  confReg_290 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  confReg_291 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  confReg_292 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  confReg_293 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  confReg_294 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  confReg_295 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  confReg_296 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  confReg_297 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  confReg_298 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  confReg_299 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  confReg_300 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  confReg_301 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  confReg_302 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  confReg_303 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  confReg_304 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  confReg_305 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  confReg_306 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  confReg_307 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  confReg_308 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  confReg_309 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  confReg_310 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  confReg_311 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  confReg_312 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  confReg_313 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  confReg_314 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  confReg_315 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  confReg_316 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  confReg_317 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  confReg_318 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  confReg_319 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  confReg_320 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  confReg_321 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  confReg_322 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  confReg_323 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  confReg_324 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  confReg_325 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  confReg_326 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  confReg_327 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  confReg_328 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  confReg_329 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  confReg_330 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  confReg_331 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  confReg_332 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  confReg_333 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  confReg_334 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  confReg_335 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  confReg_336 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  confReg_337 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  confReg_338 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  confReg_339 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  confReg_340 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  confReg_341 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  confReg_342 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  confReg_343 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  confReg_344 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  confReg_345 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  confReg_346 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  confReg_347 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  confReg_348 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  confReg_349 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  confReg_350 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  confReg_351 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  confReg_352 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  confReg_353 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  confReg_354 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  confReg_355 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  confReg_356 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  confReg_357 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  confReg_358 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  confReg_359 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  confReg_360 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  confReg_361 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  confReg_362 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  confReg_363 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  confReg_364 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  confReg_365 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  confReg_366 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  confReg_367 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  confReg_368 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  confReg_369 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  confReg_370 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  confReg_371 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  confReg_372 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  confReg_373 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  confReg_374 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  confReg_375 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  confReg_376 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  confReg_377 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  confReg_378 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  confReg_379 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  confReg_380 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  confReg_381 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  confReg_382 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  confReg_383 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  confReg_384 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  confReg_385 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  confReg_386 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  confReg_387 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  confReg_388 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  confReg_389 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  confReg_390 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  confReg_391 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  confReg_392 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  confReg_393 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  confReg_394 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  confReg_395 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  confReg_396 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  confReg_397 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  confReg_398 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  confReg_399 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  confReg_400 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  confReg_401 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  confReg_402 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  confReg_403 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  confReg_404 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  confReg_405 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  confReg_406 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  confReg_407 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  confReg_408 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  confReg_409 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  confReg_410 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  confReg_411 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  confReg_412 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  confReg_413 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  confReg_414 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  confReg_415 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  confReg_416 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  confReg_417 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  confReg_418 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  confReg_419 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  confReg_420 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  confReg_421 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  confReg_422 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  confReg_423 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  confReg_424 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  confReg_425 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  confReg_426 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  confReg_427 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  confReg_428 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  confReg_429 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  confReg_430 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  confReg_431 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  confReg_432 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  confReg_433 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  confReg_434 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  confReg_435 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  confReg_436 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  confReg_437 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  confReg_438 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  confReg_439 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  confReg_440 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  confReg_441 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  confReg_442 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  confReg_443 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  confReg_444 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  confReg_445 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  confReg_446 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  confReg_447 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  confReg_448 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  confReg_449 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  confReg_450 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  confReg_451 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  confReg_452 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  confReg_453 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  confReg_454 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  confReg_455 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  confReg_456 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  confReg_457 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  confReg_458 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  confReg_459 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  confReg_460 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  confReg_461 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  confReg_462 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  confReg_463 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  confReg_464 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  confReg_465 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  confReg_466 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  confReg_467 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  confReg_468 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  confReg_469 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  confReg_470 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  confReg_471 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  confReg_472 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  confReg_473 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  confReg_474 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  confReg_475 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  confReg_476 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  confReg_477 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  confReg_478 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  confReg_479 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  confReg_480 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  confReg_481 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  confReg_482 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  confReg_483 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  confReg_484 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  confReg_485 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  confReg_486 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  confReg_487 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  confReg_488 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  confReg_489 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  confReg_490 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  confReg_491 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  confReg_492 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  confReg_493 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  confReg_494 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  confReg_495 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  confReg_496 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  confReg_497 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  confReg_498 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  confReg_499 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  confReg_500 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  confReg_501 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  confReg_502 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  confReg_503 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  confReg_504 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  confReg_505 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  confReg_506 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  confReg_507 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  confReg_508 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  confReg_509 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  confReg_510 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  confReg_511 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  confReg_512 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  confReg_513 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  confReg_514 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  confReg_515 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  confReg_516 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  confReg_517 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  confReg_518 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  confReg_519 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  confReg_520 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  confReg_521 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  confReg_522 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  confReg_523 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  confReg_524 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  confReg_525 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  confReg_526 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  confReg_527 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  confReg_528 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  confReg_529 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  confReg_530 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  confReg_531 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  confReg_532 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  confReg_533 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  confReg_534 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  confReg_535 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  confReg_536 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  confReg_537 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  confReg_538 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  confReg_539 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  confReg_540 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  confReg_541 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  confReg_542 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  confReg_543 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  confReg_544 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  confReg_545 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  confReg_546 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  confReg_547 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  confReg_548 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  confReg_549 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  confReg_550 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  confReg_551 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  confReg_552 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  confReg_553 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  confReg_554 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  confReg_555 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  confReg_556 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  confReg_557 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  confReg_558 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  confReg_559 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  confReg_560 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  confReg_561 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  confReg_562 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  confReg_563 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  confReg_564 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  confReg_565 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  confReg_566 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  confReg_567 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  confReg_568 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  confReg_569 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  confReg_570 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  confReg_571 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  confReg_572 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  confReg_573 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  confReg_574 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  confReg_575 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  confReg_576 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  confReg_577 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  confReg_578 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  confReg_579 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  confReg_580 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  confReg_581 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  confReg_582 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  confReg_583 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  confReg_584 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  confReg_585 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  confReg_586 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  confReg_587 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  confReg_588 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  confReg_589 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  confReg_590 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  confReg_591 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  confReg_592 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  confReg_593 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  confReg_594 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  confReg_595 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  confReg_596 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  confReg_597 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  confReg_598 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  confReg_599 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  confReg_600 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  confReg_601 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  confReg_602 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  confReg_603 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  confReg_604 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  confReg_605 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  confReg_606 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  confReg_607 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  confReg_608 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  confReg_609 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  confReg_610 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  confReg_611 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  confReg_612 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  confReg_613 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  confReg_614 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  confReg_615 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  confReg_616 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  confReg_617 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  confReg_618 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  confReg_619 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  confReg_620 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  confReg_621 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  confReg_622 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  confReg_623 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  confReg_624 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  confReg_625 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  confReg_626 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  confReg_627 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  confReg_628 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  confReg_629 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  confReg_630 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  confReg_631 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  confReg_632 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  confReg_633 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  confReg_634 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  confReg_635 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  confReg_636 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  confReg_637 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  confReg_638 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  confReg_639 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  confReg_640 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  confReg_641 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  confReg_642 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  confReg_643 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  confReg_644 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  confReg_645 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  confReg_646 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  confReg_647 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  confReg_648 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  confReg_649 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  confReg_650 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  confReg_651 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  confReg_652 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  confReg_653 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  confReg_654 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  confReg_655 = _RAND_655[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MuxNInput_28_SCAOptCB(
  input  [27:0] io_in,
  input  [4:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [31:0] OPinMux_in; // @[MuxListTest.scala 44:28]
  wire [4:0] OPinMux_sel; // @[MuxListTest.scala 44:28]
  wire  OPinMux_o; // @[MuxListTest.scala 44:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux32C OPinMux ( // @[MuxListTest.scala 44:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{4'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_24_SCAOptCB(
  input  [23:0] io_in,
  input  [4:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [31:0] OPinMux_in; // @[MuxListTest.scala 44:28]
  wire [4:0] OPinMux_sel; // @[MuxListTest.scala 44:28]
  wire  OPinMux_o; // @[MuxListTest.scala 44:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux32C OPinMux ( // @[MuxListTest.scala 44:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{8'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_22_SCAOptCB(
  input  [21:0] io_in,
  input  [4:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [31:0] OPinMux_in; // @[MuxListTest.scala 44:28]
  wire [4:0] OPinMux_sel; // @[MuxListTest.scala 44:28]
  wire  OPinMux_o; // @[MuxListTest.scala 44:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux32C OPinMux ( // @[MuxListTest.scala 44:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{10'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_26_SCAOptCB(
  input  [25:0] io_in,
  input  [4:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_cnstClk,
  input         io_arst
);
  wire [31:0] OPinMux_in; // @[MuxListTest.scala 44:28]
  wire [4:0] OPinMux_sel; // @[MuxListTest.scala 44:28]
  wire  OPinMux_o; // @[MuxListTest.scala 44:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux32C OPinMux ( // @[MuxListTest.scala 44:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{6'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_1_SCAOptCB(
  input   io_in,
  input   io_config,
  output  io_out,
  input   io_loopBreak,
  input   io_cnstClk,
  input   io_arst
);
  wire [1:0] OPinMux_in; // @[MuxListTest.scala 40:28]
  wire  OPinMux_sel; // @[MuxListTest.scala 40:28]
  wire  OPinMux_o; // @[MuxListTest.scala 40:28]
  wire  lbCBFlop_d; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_rb; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_clk; // @[MuxListTest.scala 59:24]
  wire  lbCBFlop_o; // @[MuxListTest.scala 59:24]
  wire  lbNor_a; // @[MuxListTest.scala 64:23]
  wire  lbNor_b; // @[MuxListTest.scala 64:23]
  wire  lbNor_o1; // @[MuxListTest.scala 64:23]
  Mux2C OPinMux ( // @[MuxListTest.scala 40:28]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  b0mfqn003hn1n02x5 lbCBFlop ( // @[MuxListTest.scala 59:24]
    .d(lbCBFlop_d),
    .rb(lbCBFlop_rb),
    .clk(lbCBFlop_clk),
    .o(lbCBFlop_o)
  );
  b0mnor002an1n04x5 lbNor ( // @[MuxListTest.scala 64:23]
    .a(lbNor_a),
    .b(lbNor_b),
    .o1(lbNor_o1)
  );
  assign io_out = ~(lbCBFlop_o | lbNor_o1); // @[MuxListTest.scala 71:15]
  assign OPinMux_in = {{1'd0}, io_in}; // @[MuxListTest.scala 53:20]
  assign OPinMux_sel = io_config; // @[MuxListTest.scala 52:21]
  assign lbCBFlop_d = OPinMux_o; // @[MuxListTest.scala 60:17]
  assign lbCBFlop_rb = io_arst; // @[MuxListTest.scala 62:18]
  assign lbCBFlop_clk = io_cnstClk; // @[MuxListTest.scala 61:19]
  assign lbNor_a = io_loopBreak; // @[MuxListTest.scala 65:16]
  assign lbNor_b = OPinMux_o; // @[MuxListTest.scala 66:16]
endmodule
module MuxNInput_O3_C6_SCAOptSB(
  input  [8:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{5'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in[8:3]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O3_C7_SCAOptSB(
  input  [9:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{5'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{1'd0}, io_in[9:3]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O3_C5_SCAOptSB(
  input  [7:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{5'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in[7:3]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O2_C5_SCAOptSB(
  input  [6:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{6'd0}, io_in[1:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in[6:2]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O0_C1_SCAOptSB(
  input        io_in,
  input  [1:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [1:0] OPinMux_in; // @[MuxListTest.scala 108:26]
  wire  OPinMux_sel; // @[MuxListTest.scala 108:26]
  wire  OPinMux_o; // @[MuxListTest.scala 108:26]
  wire [1:0] chanMux_in; // @[MuxListTest.scala 129:26]
  wire  chanMux_sel; // @[MuxListTest.scala 129:26]
  wire  chanMux_o; // @[MuxListTest.scala 129:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux2C OPinMux ( // @[MuxListTest.scala 108:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux2C chanMux ( // @[MuxListTest.scala 129:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = 2'h0; // @[MuxListTest.scala 125:22]
  assign OPinMux_sel = io_config[0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{1'd0}, io_in}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[1] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O2_C6_SCAOptSB(
  input  [7:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{6'd0}, io_in[1:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in[7:2]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O4_C6_SCAOptSB(
  input  [9:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{4'd0}, io_in[3:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{2'd0}, io_in[9:4]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O4_C7_SCAOptSB(
  input  [10:0] io_in,
  input  [3:0]  io_config,
  output        io_out,
  input         io_loopBreak,
  input         io_ioGndBle,
  input         io_cnstClk,
  input         io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{4'd0}, io_in[3:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{1'd0}, io_in[10:4]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O3_C4_SCAOptSB(
  input  [6:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{1'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = io_in[6:3]; // @[MuxListTest.scala 145:30]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O4_C5_SCAOptSB(
  input  [8:0] io_in,
  input  [3:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [7:0] OPinMux_in; // @[MuxListTest.scala 110:26]
  wire [2:0] OPinMux_sel; // @[MuxListTest.scala 110:26]
  wire  OPinMux_o; // @[MuxListTest.scala 110:26]
  wire [7:0] chanMux_in; // @[MuxListTest.scala 131:26]
  wire [2:0] chanMux_sel; // @[MuxListTest.scala 131:26]
  wire  chanMux_o; // @[MuxListTest.scala 131:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux8C OPinMux ( // @[MuxListTest.scala 110:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux8C chanMux ( // @[MuxListTest.scala 131:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{4'd0}, io_in[3:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[2:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in[8:4]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[2:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[3] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O4_C1_SCAOptSB(
  input  [4:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = io_in[3:0]; // @[MuxListTest.scala 123:30]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in[4]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module MuxNInput_O3_C1_SCAOptSB(
  input  [3:0] io_in,
  input  [2:0] io_config,
  output       io_out,
  input        io_loopBreak,
  input        io_ioGndBle,
  input        io_cnstClk,
  input        io_arst
);
  wire [3:0] OPinMux_in; // @[MuxListTest.scala 109:26]
  wire [1:0] OPinMux_sel; // @[MuxListTest.scala 109:26]
  wire  OPinMux_o; // @[MuxListTest.scala 109:26]
  wire [3:0] chanMux_in; // @[MuxListTest.scala 130:26]
  wire [1:0] chanMux_sel; // @[MuxListTest.scala 130:26]
  wire  chanMux_o; // @[MuxListTest.scala 130:26]
  wire  lbCBMux_a; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_b; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_sa; // @[MuxListTest.scala 151:22]
  wire  lbCBMux_o; // @[MuxListTest.scala 151:22]
  wire  lbSBFlop_d; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_rb; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_clk; // @[MuxListTest.scala 152:22]
  wire  lbSBFlop_o; // @[MuxListTest.scala 152:22]
  Mux4C OPinMux ( // @[MuxListTest.scala 109:26]
    .in(OPinMux_in),
    .sel(OPinMux_sel),
    .o(OPinMux_o)
  );
  Mux4C chanMux ( // @[MuxListTest.scala 130:26]
    .in(chanMux_in),
    .sel(chanMux_sel),
    .o(chanMux_o)
  );
  b0mmbn022ah1n02x5 lbCBMux ( // @[MuxListTest.scala 151:22]
    .a(lbCBMux_a),
    .b(lbCBMux_b),
    .sa(lbCBMux_sa),
    .o(lbCBMux_o)
  );
  b0mfqn003hn1n02x5 lbSBFlop ( // @[MuxListTest.scala 152:22]
    .d(lbSBFlop_d),
    .rb(lbSBFlop_rb),
    .clk(lbSBFlop_clk),
    .o(lbSBFlop_o)
  );
  assign io_out = lbCBMux_o | lbSBFlop_o & io_ioGndBle; // @[MuxListTest.scala 160:25]
  assign OPinMux_in = {{1'd0}, io_in[2:0]}; // @[MuxListTest.scala 123:22]
  assign OPinMux_sel = io_config[1:0]; // @[MuxListTest.scala 121:33]
  assign chanMux_in = {{3'd0}, io_in[3]}; // @[MuxListTest.scala 145:22]
  assign chanMux_sel = io_config[1:0]; // @[MuxListTest.scala 143:33]
  assign lbCBMux_a = OPinMux_o; // @[MuxListTest.scala 158:15]
  assign lbCBMux_b = chanMux_o; // @[MuxListTest.scala 159:15]
  assign lbCBMux_sa = io_config[2] | io_loopBreak; // @[MuxListTest.scala 157:43]
  assign lbSBFlop_d = ~(chanMux_o & OPinMux_o); // @[MuxListTest.scala 153:18]
  assign lbSBFlop_rb = io_arst; // @[MuxListTest.scala 155:16]
  assign lbSBFlop_clk = io_cnstClk; // @[MuxListTest.scala 154:17]
endmodule
module Tile_7_1_clbmultile(
  input          clock,
  input          reset,
  input          IN_OPIN_N15079_73,
  input          IN_OPIN_N15080_74,
  input          IN_OPIN_N15081_75,
  input          IN_OPIN_N15082_76,
  input          IN_OPIN_N15083_77,
  input          IN_OPIN_N15084_78,
  input          IN_OPIN_N15085_79,
  input          IN_OPIN_N15086_80,
  input          IN_OPIN_N15095_89,
  input          IN_OPIN_N15096_90,
  input          IN_OPIN_N15097_91,
  input          IN_OPIN_N15098_92,
  input          IN_OPIN_N15099_93,
  input          IN_OPIN_N15100_94,
  input          IN_OPIN_N15101_95,
  input          IN_OPIN_N15102_96,
  input          IN_OPIN_N15103_97,
  input          IN_OPIN_N15104_98,
  input          IN_OPIN_N15105_99,
  input          IN_OPIN_N15106_100,
  input          IN_OPIN_N15107_101,
  input          IN_OPIN_N15108_102,
  input          IN_OPIN_N15109_103,
  input          IN_OPIN_N15110_104,
  input          IN_OPIN_N15111_105,
  input          IN_OPIN_N15112_106,
  input          IN_OPIN_N15113_107,
  input          IN_OPIN_N15114_108,
  input          IN_OPIN_N15115_109,
  input          IN_OPIN_N15116_110,
  input          IN_OPIN_N15117_111,
  input          IN_OPIN_N15118_112,
  input          IN_OPIN_N15119_113,
  input          IN_OPIN_N15120_114,
  input          IN_OPIN_N15121_115,
  input          IN_OPIN_N15122_116,
  input          IN_OPIN_N15123_117,
  input          IN_OPIN_N15124_118,
  input          IN_OPIN_N15125_119,
  input          IN_OPIN_N15126_120,
  input          IN_OPIN_N17283_81,
  input          IN_OPIN_N17284_82,
  input          IN_OPIN_N17285_83,
  input          IN_OPIN_N17286_84,
  input          IN_OPIN_N17287_85,
  input          IN_OPIN_N17288_86,
  input          IN_OPIN_N17289_87,
  input          IN_OPIN_N17290_88,
  input          IN_CHANX_N23682_0,
  input          IN_CHANX_N23684_8,
  input          IN_CHANX_N23686_16,
  input          IN_CHANX_N23688_24,
  input          IN_CHANX_N23690_32,
  input          IN_CHANX_N23692_40,
  input          IN_CHANX_N23694_48,
  input          IN_CHANX_N23696_56,
  input          IN_CHANX_N23698_64,
  input          IN_CHANX_N23700_72,
  input          IN_CHANX_N23702_80,
  input          IN_CHANX_N23704_88,
  input          IN_CHANX_N23706_96,
  input          IN_CHANX_N23712_2,
  input          IN_CHANX_N23713_3,
  input          IN_CHANX_N23714_10,
  input          IN_CHANX_N23715_11,
  input          IN_CHANX_N23716_18,
  input          IN_CHANX_N23717_19,
  input          IN_CHANX_N23718_26,
  input          IN_CHANX_N23719_27,
  input          IN_CHANX_N23720_34,
  input          IN_CHANX_N23721_35,
  input          IN_CHANX_N23722_42,
  input          IN_CHANX_N23723_43,
  input          IN_CHANX_N23724_50,
  input          IN_CHANX_N23725_51,
  input          IN_CHANX_N23726_58,
  input          IN_CHANX_N23727_59,
  input          IN_CHANX_N23728_66,
  input          IN_CHANX_N23729_67,
  input          IN_CHANX_N23730_74,
  input          IN_CHANX_N23731_75,
  input          IN_CHANX_N23732_82,
  input          IN_CHANX_N23733_83,
  input          IN_CHANX_N23742_4,
  input          IN_CHANX_N23743_5,
  input          IN_CHANX_N23744_12,
  input          IN_CHANX_N23745_13,
  input          IN_CHANX_N23746_20,
  input          IN_CHANX_N23747_21,
  input          IN_CHANX_N23748_28,
  input          IN_CHANX_N23749_29,
  input          IN_CHANX_N23750_36,
  input          IN_CHANX_N23751_37,
  input          IN_CHANX_N23752_44,
  input          IN_CHANX_N23753_45,
  input          IN_CHANX_N23754_52,
  input          IN_CHANX_N23755_53,
  input          IN_CHANX_N23756_60,
  input          IN_CHANX_N23757_61,
  input          IN_CHANX_N23758_68,
  input          IN_CHANX_N23759_69,
  input          IN_CHANX_N23760_76,
  input          IN_CHANX_N23761_77,
  input          IN_CHANX_N23766_100,
  input          IN_CHANX_N23768_104,
  input          IN_CHANX_N23770_6,
  input          IN_CHANX_N23771_7,
  input          IN_CHANX_N23772_14,
  input          IN_CHANX_N23773_15,
  input          IN_CHANX_N23774_22,
  input          IN_CHANX_N23775_23,
  input          IN_CHANX_N23776_30,
  input          IN_CHANX_N23777_31,
  input          IN_CHANX_N23778_38,
  input          IN_CHANX_N23779_39,
  input          IN_CHANX_N23780_46,
  input          IN_CHANX_N23781_47,
  input          IN_CHANX_N23782_54,
  input          IN_CHANX_N23783_55,
  input          IN_CHANX_N23784_62,
  input          IN_CHANX_N23785_63,
  input          IN_CHANX_N23786_70,
  input          IN_CHANX_N23787_71,
  input          IN_CHANX_N23788_78,
  input          IN_CHANX_N23789_79,
  input          IN_CHANX_N23790_86,
  input          IN_CHANX_N23791_87,
  input          IN_CHANX_N23792_94,
  input          IN_CHANX_N23793_95,
  input          IN_CHANX_N23794_102,
  input          IN_CHANX_N23795_103,
  input          IN_CHANX_N23796_106,
  input          IN_CHANX_N23797_107,
  input          IN_CHANX_N23799_1,
  input          IN_CHANX_N23801_9,
  input          IN_CHANX_N23803_17,
  input          IN_CHANX_N23809_41,
  input          IN_CHANX_N23813_57,
  input          IN_CHANX_N23821_89,
  input          IN_CHANX_N23823_97,
  input          IN_CHANX_N23825_101,
  input          IN_CHANX_N23827_105,
  input          IN_CHANY_N30078_0,
  input          IN_CHANY_N30080_2,
  input          IN_CHANY_N30081_3,
  input          IN_CHANY_N30082_4,
  input          IN_CHANY_N30083_5,
  input          IN_CHANY_N30084_6,
  input          IN_CHANY_N30085_7,
  input          IN_CHANY_N30086_8,
  input          IN_CHANY_N30088_10,
  input          IN_CHANY_N30089_11,
  input          IN_CHANY_N30090_12,
  input          IN_CHANY_N30091_13,
  input          IN_CHANY_N30092_14,
  input          IN_CHANY_N30093_15,
  input          IN_CHANY_N30094_16,
  input          IN_CHANY_N30096_18,
  input          IN_CHANY_N30097_19,
  input          IN_CHANY_N30098_20,
  input          IN_CHANY_N30099_21,
  input          IN_CHANY_N30100_22,
  input          IN_CHANY_N30101_23,
  input          IN_CHANY_N30102_24,
  input          IN_CHANY_N30104_26,
  input          IN_CHANY_N30105_27,
  input          IN_CHANY_N30106_28,
  input          IN_CHANY_N30107_29,
  input          IN_CHANY_N30108_30,
  input          IN_CHANY_N30109_31,
  input          IN_CHANY_N30110_32,
  input          IN_CHANY_N30112_34,
  input          IN_CHANY_N30113_35,
  input          IN_CHANY_N30114_36,
  input          IN_CHANY_N30115_37,
  input          IN_CHANY_N30116_38,
  input          IN_CHANY_N30117_39,
  input          IN_CHANY_N30118_40,
  input          IN_CHANY_N30120_42,
  input          IN_CHANY_N30121_43,
  input          IN_CHANY_N30122_44,
  input          IN_CHANY_N30123_45,
  input          IN_CHANY_N30124_46,
  input          IN_CHANY_N30125_47,
  input          IN_CHANY_N30126_48,
  input          IN_CHANY_N30128_50,
  input          IN_CHANY_N30129_51,
  input          IN_CHANY_N30130_52,
  input          IN_CHANY_N30131_53,
  input          IN_CHANY_N30132_54,
  input          IN_CHANY_N30133_55,
  input          IN_CHANY_N30134_56,
  input          IN_CHANY_N30136_58,
  input          IN_CHANY_N30137_59,
  input          IN_CHANY_N30138_60,
  input          IN_CHANY_N30139_61,
  input          IN_CHANY_N30140_62,
  input          IN_CHANY_N30141_63,
  input          IN_CHANY_N30142_64,
  input          IN_CHANY_N30144_66,
  input          IN_CHANY_N30145_67,
  input          IN_CHANY_N30146_68,
  input          IN_CHANY_N30147_69,
  input          IN_CHANY_N30148_70,
  input          IN_CHANY_N30149_71,
  input          IN_CHANY_N30150_72,
  input          IN_CHANY_N30152_74,
  input          IN_CHANY_N30153_75,
  input          IN_CHANY_N30154_76,
  input          IN_CHANY_N30155_77,
  input          IN_CHANY_N30156_78,
  input          IN_CHANY_N30157_79,
  input          IN_CHANY_N30158_80,
  input          IN_CHANY_N30160_82,
  input          IN_CHANY_N30161_83,
  input          IN_CHANY_N30162_84,
  input          IN_CHANY_N30163_85,
  input          IN_CHANY_N30164_86,
  input          IN_CHANY_N30165_87,
  input          IN_CHANY_N30166_88,
  input          IN_CHANY_N30168_90,
  input          IN_CHANY_N30169_91,
  input          IN_CHANY_N30170_92,
  input          IN_CHANY_N30171_93,
  input          IN_CHANY_N30172_94,
  input          IN_CHANY_N30173_95,
  input          IN_CHANY_N30174_96,
  input          IN_CHANY_N30176_98,
  input          IN_CHANY_N30177_99,
  input          IN_CHANY_N30178_100,
  input          IN_CHANY_N30180_102,
  input          IN_CHANY_N30181_103,
  input          IN_CHANY_N30182_104,
  input          IN_CHANY_N30184_106,
  input          IN_CHANY_N30185_107,
  input          IN_CHANY_N30193_25,
  input          IN_CHANY_N30195_33,
  input          IN_CHANY_N30199_49,
  input          IN_CHANY_N30201_57,
  input          IN_CHANY_N30205_73,
  input          IN_CHANY_N30209_89,
  input          IN_CHANY_N30211_97,
  input          IN_CHANY_N30213_101,
  input          IN_CHANY_N30215_105,
  output         OUT_CHANX_N23695_49,
  output         OUT_OPIN_N14842_80,
  output         OUT_CHANX_N23824_100,
  output         OUT_OPIN_N14846_84,
  output         OUT_OPIN_N14850_88,
  output         OUT_CHANY_N30196_40,
  output         OUT_CHANX_N23802_16,
  output         OUT_CHANX_N23691_33,
  output         OUT_OPIN_N14847_85,
  output         OUT_CHANY_N30175_97,
  output         OUT_CHANY_N30212_100,
  output         OUT_CHANX_N23798_0,
  output         OUT_CHANY_N30198_48,
  output         OUT_OPIN_N14840_78,
  output         OUT_CHANX_N23685_9,
  output         OUT_OPIN_N14844_82,
  output         OUT_CHANX_N23816_72,
  output         OUT_CHANX_N23769_105,
  output         OUT_CHANX_N23683_1,
  output         OUT_CHANX_N23826_104,
  output         OUT_CHANX_N23810_48,
  output         OUT_OPIN_N14837_75,
  output         OUT_CHANX_N23822_96,
  output         OUT_CHANY_N30204_72,
  output         OUT_OPIN_N14836_74,
  output         OUT_CHANX_N23800_8,
  output         OUT_CHANX_N23804_24,
  output         OUT_CHANX_N23812_56,
  output         OUT_OPIN_N14845_83,
  output         OUT_CHANY_N30190_16,
  output         OUT_CHANY_N30159_81,
  output         OUT_CHANY_N30214_104,
  output         OUT_CHANX_N23707_97,
  output         OUT_OPIN_N14843_81,
  output         OUT_CHANX_N23808_40,
  output         OUT_CHANY_N30087_9,
  output         OUT_CHANY_N30206_80,
  output         OUT_CHANY_N30208_88,
  output         OUT_CHANY_N30119_41,
  output         OUT_OPIN_N14849_87,
  output         OUT_CHANY_N30192_24,
  output         OUT_CHANY_N30143_65,
  output         OUT_CHANY_N30095_17,
  output         OUT_CHANY_N30186_0,
  output         OUT_OPIN_N14835_73,
  output         OUT_CHANX_N23701_73,
  output         OUT_CHANX_N23689_25,
  output         OUT_CHANX_N23814_64,
  output         OUT_CHANX_N23697_57,
  output         OUT_CHANX_N23687_17,
  output         OUT_CHANY_N30202_64,
  output         OUT_OPIN_N14841_79,
  output         OUT_OPIN_N14838_76,
  output         OUT_CHANX_N23699_65,
  output         OUT_CHANX_N23767_101,
  output         OUT_CHANY_N30194_32,
  output         OUT_CHANY_N30188_8,
  output         OUT_CHANX_N23818_80,
  output         OUT_CHANY_N30210_96,
  output         OUT_OPIN_N14839_77,
  output         OUT_CHANX_N23703_81,
  output         OUT_CHANY_N30200_56,
  output         OUT_CHANY_N30167_89,
  output         OUT_OPIN_N14848_86,
  output         OUT_CHANX_N23693_41,
  output         OUT_CHANX_N23820_88,
  output         OUT_CHANX_N23806_32,
  output         OUT_CHANY_N30183_105,
  output         OUT_CHANX_N23705_89,
  output         OUT_CHANY_N30179_101,
  output [652:0] ioConf_confOut,
  input  [15:0]  ioConf_scan_in,
  input          ioConf_scan_en,
  output [15:0]  ioConf_scan_out,
  input          ctrlSignals_gndBlkOuts,
  input          ctrlSignals_loopBreak,
  input          ctrlSignals_arst,
  input          ctrlSignals_confClock,
  input          ctrlSignals_constClock
);
  wire  logicBlock_IPIN_0; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_1; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_2; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_3; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_4; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_5; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_6; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_7; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_8; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_9; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_10; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_11; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_12; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_13; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_14; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_15; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_16; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_17; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_18; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_19; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_20; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_21; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_22; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_23; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_24; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_25; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_26; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_27; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_28; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_29; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_30; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_31; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_32; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_33; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_34; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_35; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_36; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_37; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_38; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_39; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_40; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_41; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_42; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_43; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_44; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_45; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_46; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_47; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_48; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_49; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_50; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_51; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_52; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_53; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_54; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_55; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_56; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_57; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_58; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_59; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_60; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_61; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_62; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_63; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_64; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_65; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_66; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_67; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_68; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_69; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_70; // @[TileFull.scala 47:37]
  wire  logicBlock_IPIN_71; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_73; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_74; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_75; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_76; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_77; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_78; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_79; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_80; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_81; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_82; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_83; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_84; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_85; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_86; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_87; // @[TileFull.scala 47:37]
  wire  logicBlock_OPIN_88; // @[TileFull.scala 47:37]
  wire  logicBlock_clock; // @[TileFull.scala 47:37]
  wire  logicBlock_reset; // @[TileFull.scala 47:37]
  wire [193:0] logicBlock_configBits; // @[TileFull.scala 47:37]
  wire  logicBlock_loopBreak; // @[TileFull.scala 47:37]
  wire  logicBlock_gndLBouts; // @[TileFull.scala 47:37]
  wire  configBlock_clock; // @[TileFull.scala 66:31]
  wire [655:0] configBlock_ioBundle_confOut; // @[TileFull.scala 66:31]
  wire [15:0] configBlock_ioBundle_scan_in; // @[TileFull.scala 66:31]
  wire  configBlock_ioBundle_scan_en; // @[TileFull.scala 66:31]
  wire [15:0] configBlock_ioBundle_scan_out; // @[TileFull.scala 66:31]
  wire [27:0] CBMux_IPIN0_N14762_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN0_N14762_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN0_N14762_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN0_N14762_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN0_N14762_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN0_N14762_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN1_N14763_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN1_N14763_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN1_N14763_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN1_N14763_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN1_N14763_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN1_N14763_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN2_N14764_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN2_N14764_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN2_N14764_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN2_N14764_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN2_N14764_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN2_N14764_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN3_N14765_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN3_N14765_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN3_N14765_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN3_N14765_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN3_N14765_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN3_N14765_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN4_N14766_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN4_N14766_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN4_N14766_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN4_N14766_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN4_N14766_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN4_N14766_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN5_N14767_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN5_N14767_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN5_N14767_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN5_N14767_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN5_N14767_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN5_N14767_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN6_N14768_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN6_N14768_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN6_N14768_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN6_N14768_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN6_N14768_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN6_N14768_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN7_N14769_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN7_N14769_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN7_N14769_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN7_N14769_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN7_N14769_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN7_N14769_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN8_N14770_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN8_N14770_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN8_N14770_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN8_N14770_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN8_N14770_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN8_N14770_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN9_N14771_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN9_N14771_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN9_N14771_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN9_N14771_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN9_N14771_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN9_N14771_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN10_N14772_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN10_N14772_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN10_N14772_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN10_N14772_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN10_N14772_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN10_N14772_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN11_N14773_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN11_N14773_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN11_N14773_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN11_N14773_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN11_N14773_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN11_N14773_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN12_N14774_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN12_N14774_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN12_N14774_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN12_N14774_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN12_N14774_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN12_N14774_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN13_N14775_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN13_N14775_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN13_N14775_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN13_N14775_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN13_N14775_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN13_N14775_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN14_N14776_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN14_N14776_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN14_N14776_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN14_N14776_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN14_N14776_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN14_N14776_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN15_N14777_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN15_N14777_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN15_N14777_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN15_N14777_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN15_N14777_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN15_N14777_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN16_N14778_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN16_N14778_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN16_N14778_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN16_N14778_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN16_N14778_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN16_N14778_io_arst; // @[TileFull.scala 102:29]
  wire [27:0] CBMux_IPIN17_N14779_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN17_N14779_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN17_N14779_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN17_N14779_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN17_N14779_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN17_N14779_io_arst; // @[TileFull.scala 102:29]
  wire [23:0] CBMux_IPIN18_N14780_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN18_N14780_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN18_N14780_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN18_N14780_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN18_N14780_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN18_N14780_io_arst; // @[TileFull.scala 102:29]
  wire [23:0] CBMux_IPIN19_N14781_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN19_N14781_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN19_N14781_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN19_N14781_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN19_N14781_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN19_N14781_io_arst; // @[TileFull.scala 102:29]
  wire [21:0] CBMux_IPIN20_N14782_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN20_N14782_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN20_N14782_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN20_N14782_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN20_N14782_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN20_N14782_io_arst; // @[TileFull.scala 102:29]
  wire [25:0] CBMux_IPIN21_N14783_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN21_N14783_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN21_N14783_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN21_N14783_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN21_N14783_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN21_N14783_io_arst; // @[TileFull.scala 102:29]
  wire [25:0] CBMux_IPIN22_N14784_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN22_N14784_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN22_N14784_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN22_N14784_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN22_N14784_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN22_N14784_io_arst; // @[TileFull.scala 102:29]
  wire [21:0] CBMux_IPIN23_N14785_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN23_N14785_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN23_N14785_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN23_N14785_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN23_N14785_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN23_N14785_io_arst; // @[TileFull.scala 102:29]
  wire [21:0] CBMux_IPIN24_N14786_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN24_N14786_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN24_N14786_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN24_N14786_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN24_N14786_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN24_N14786_io_arst; // @[TileFull.scala 102:29]
  wire [21:0] CBMux_IPIN25_N14787_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN25_N14787_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN25_N14787_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN25_N14787_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN25_N14787_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN25_N14787_io_arst; // @[TileFull.scala 102:29]
  wire [25:0] CBMux_IPIN26_N14788_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN26_N14788_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN26_N14788_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN26_N14788_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN26_N14788_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN26_N14788_io_arst; // @[TileFull.scala 102:29]
  wire [25:0] CBMux_IPIN27_N14789_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN27_N14789_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN27_N14789_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN27_N14789_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN27_N14789_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN27_N14789_io_arst; // @[TileFull.scala 102:29]
  wire [25:0] CBMux_IPIN28_N14790_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN28_N14790_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN28_N14790_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN28_N14790_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN28_N14790_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN28_N14790_io_arst; // @[TileFull.scala 102:29]
  wire [21:0] CBMux_IPIN29_N14791_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN29_N14791_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN29_N14791_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN29_N14791_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN29_N14791_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN29_N14791_io_arst; // @[TileFull.scala 102:29]
  wire [21:0] CBMux_IPIN30_N14792_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN30_N14792_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN30_N14792_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN30_N14792_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN30_N14792_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN30_N14792_io_arst; // @[TileFull.scala 102:29]
  wire [25:0] CBMux_IPIN31_N14793_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN31_N14793_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN31_N14793_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN31_N14793_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN31_N14793_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN31_N14793_io_arst; // @[TileFull.scala 102:29]
  wire [25:0] CBMux_IPIN32_N14794_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN32_N14794_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN32_N14794_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN32_N14794_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN32_N14794_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN32_N14794_io_arst; // @[TileFull.scala 102:29]
  wire [25:0] CBMux_IPIN33_N14795_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN33_N14795_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN33_N14795_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN33_N14795_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN33_N14795_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN33_N14795_io_arst; // @[TileFull.scala 102:29]
  wire [21:0] CBMux_IPIN34_N14796_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN34_N14796_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN34_N14796_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN34_N14796_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN34_N14796_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN34_N14796_io_arst; // @[TileFull.scala 102:29]
  wire [21:0] CBMux_IPIN35_N14797_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN35_N14797_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN35_N14797_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN35_N14797_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN35_N14797_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN35_N14797_io_arst; // @[TileFull.scala 102:29]
  wire [21:0] CBMux_IPIN36_N14798_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN36_N14798_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN36_N14798_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN36_N14798_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN36_N14798_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN36_N14798_io_arst; // @[TileFull.scala 102:29]
  wire [25:0] CBMux_IPIN37_N14799_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN37_N14799_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN37_N14799_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN37_N14799_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN37_N14799_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN37_N14799_io_arst; // @[TileFull.scala 102:29]
  wire [25:0] CBMux_IPIN38_N14800_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN38_N14800_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN38_N14800_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN38_N14800_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN38_N14800_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN38_N14800_io_arst; // @[TileFull.scala 102:29]
  wire [21:0] CBMux_IPIN39_N14801_io_in; // @[TileFull.scala 102:29]
  wire [4:0] CBMux_IPIN39_N14801_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN39_N14801_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN39_N14801_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN39_N14801_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN39_N14801_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN40_N14802_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN40_N14802_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN40_N14802_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN40_N14802_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN40_N14802_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN40_N14802_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN41_N14803_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN41_N14803_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN41_N14803_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN41_N14803_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN41_N14803_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN41_N14803_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN42_N14804_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN42_N14804_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN42_N14804_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN42_N14804_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN42_N14804_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN42_N14804_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN43_N14805_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN43_N14805_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN43_N14805_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN43_N14805_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN43_N14805_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN43_N14805_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN44_N14806_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN44_N14806_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN44_N14806_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN44_N14806_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN44_N14806_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN44_N14806_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN45_N14807_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN45_N14807_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN45_N14807_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN45_N14807_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN45_N14807_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN45_N14807_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN46_N14808_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN46_N14808_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN46_N14808_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN46_N14808_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN46_N14808_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN46_N14808_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN47_N14809_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN47_N14809_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN47_N14809_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN47_N14809_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN47_N14809_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN47_N14809_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN48_N14810_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN48_N14810_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN48_N14810_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN48_N14810_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN48_N14810_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN48_N14810_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN49_N14811_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN49_N14811_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN49_N14811_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN49_N14811_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN49_N14811_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN49_N14811_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN50_N14812_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN50_N14812_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN50_N14812_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN50_N14812_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN50_N14812_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN50_N14812_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN51_N14813_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN51_N14813_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN51_N14813_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN51_N14813_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN51_N14813_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN51_N14813_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN52_N14814_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN52_N14814_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN52_N14814_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN52_N14814_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN52_N14814_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN52_N14814_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN53_N14815_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN53_N14815_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN53_N14815_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN53_N14815_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN53_N14815_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN53_N14815_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN54_N14816_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN54_N14816_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN54_N14816_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN54_N14816_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN54_N14816_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN54_N14816_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN55_N14817_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN55_N14817_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN55_N14817_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN55_N14817_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN55_N14817_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN55_N14817_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN56_N14818_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN56_N14818_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN56_N14818_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN56_N14818_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN56_N14818_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN56_N14818_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN57_N14819_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN57_N14819_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN57_N14819_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN57_N14819_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN57_N14819_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN57_N14819_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN58_N14820_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN58_N14820_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN58_N14820_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN58_N14820_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN58_N14820_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN58_N14820_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN59_N14821_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN59_N14821_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN59_N14821_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN59_N14821_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN59_N14821_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN59_N14821_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN60_N14822_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN60_N14822_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN60_N14822_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN60_N14822_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN60_N14822_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN60_N14822_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN61_N14823_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN61_N14823_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN61_N14823_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN61_N14823_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN61_N14823_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN61_N14823_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN62_N14824_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN62_N14824_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN62_N14824_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN62_N14824_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN62_N14824_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN62_N14824_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN63_N14825_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN63_N14825_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN63_N14825_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN63_N14825_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN63_N14825_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN63_N14825_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN64_N14826_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN64_N14826_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN64_N14826_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN64_N14826_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN64_N14826_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN64_N14826_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN65_N14827_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN65_N14827_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN65_N14827_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN65_N14827_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN65_N14827_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN65_N14827_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN66_N14828_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN66_N14828_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN66_N14828_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN66_N14828_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN66_N14828_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN66_N14828_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN67_N14829_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN67_N14829_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN67_N14829_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN67_N14829_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN67_N14829_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN67_N14829_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN68_N14830_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN68_N14830_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN68_N14830_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN68_N14830_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN68_N14830_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN68_N14830_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN69_N14831_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN69_N14831_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN69_N14831_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN69_N14831_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN69_N14831_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN69_N14831_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN70_N14832_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN70_N14832_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN70_N14832_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN70_N14832_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN70_N14832_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN70_N14832_io_arst; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN71_N14833_io_in; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN71_N14833_io_config; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN71_N14833_io_out; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN71_N14833_io_loopBreak; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN71_N14833_io_cnstClk; // @[TileFull.scala 102:29]
  wire  CBMux_IPIN71_N14833_io_arst; // @[TileFull.scala 102:29]
  wire [8:0] SBMux_C1_N23683_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C1_N23683_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C1_N23683_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C1_N23683_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C1_N23683_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C1_N23683_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C1_N23683_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [9:0] SBMux_C9_N23685_O_3_C_7_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C9_N23685_O_3_C_7_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C9_N23685_O_3_C_7_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C9_N23685_O_3_C_7_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C9_N23685_O_3_C_7_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C9_N23685_O_3_C_7_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C9_N23685_O_3_C_7_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C17_N23687_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C17_N23687_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C17_N23687_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C17_N23687_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C17_N23687_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C17_N23687_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C17_N23687_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C25_N23689_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C25_N23689_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C25_N23689_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C25_N23689_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C25_N23689_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C25_N23689_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C25_N23689_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [9:0] SBMux_C33_N23691_O_3_C_7_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C33_N23691_O_3_C_7_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C33_N23691_O_3_C_7_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C33_N23691_O_3_C_7_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C33_N23691_O_3_C_7_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C33_N23691_O_3_C_7_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C33_N23691_O_3_C_7_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C41_N23693_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C41_N23693_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C41_N23693_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C41_N23693_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C41_N23693_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C41_N23693_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C41_N23693_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [7:0] SBMux_C49_N23695_O_3_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C49_N23695_O_3_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C49_N23695_O_3_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C49_N23695_O_3_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C49_N23695_O_3_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C49_N23695_O_3_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C49_N23695_O_3_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C57_N23697_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C57_N23697_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C57_N23697_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C57_N23697_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C57_N23697_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C57_N23697_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C57_N23697_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C65_N23699_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C65_N23699_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C65_N23699_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C65_N23699_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C65_N23699_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C65_N23699_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C65_N23699_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C73_N23701_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C73_N23701_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C73_N23701_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C73_N23701_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C73_N23701_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C73_N23701_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C73_N23701_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [6:0] SBMux_C81_N23703_O_2_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C81_N23703_O_2_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C81_N23703_O_2_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C81_N23703_O_2_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C81_N23703_O_2_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C81_N23703_O_2_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C81_N23703_O_2_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [7:0] SBMux_C89_N23705_O_3_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C89_N23705_O_3_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C89_N23705_O_3_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C89_N23705_O_3_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C89_N23705_O_3_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C89_N23705_O_3_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C89_N23705_O_3_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [6:0] SBMux_C97_N23707_O_2_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C97_N23707_O_2_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C97_N23707_O_2_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C97_N23707_O_2_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C97_N23707_O_2_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C97_N23707_O_2_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C97_N23707_O_2_C_5_io_arst; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N23767_O_0_C_1_io_in; // @[TileFull.scala 141:27]
  wire [1:0] SBMux_C101_N23767_O_0_C_1_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N23767_O_0_C_1_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N23767_O_0_C_1_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N23767_O_0_C_1_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N23767_O_0_C_1_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N23767_O_0_C_1_io_arst; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N23769_O_0_C_1_io_in; // @[TileFull.scala 141:27]
  wire [1:0] SBMux_C105_N23769_O_0_C_1_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N23769_O_0_C_1_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N23769_O_0_C_1_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N23769_O_0_C_1_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N23769_O_0_C_1_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N23769_O_0_C_1_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C0_N23798_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C0_N23798_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C0_N23798_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C0_N23798_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C0_N23798_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C0_N23798_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C0_N23798_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C8_N23800_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C8_N23800_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C8_N23800_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C8_N23800_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C8_N23800_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C8_N23800_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C8_N23800_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C16_N23802_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C16_N23802_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C16_N23802_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C16_N23802_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C16_N23802_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C16_N23802_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C16_N23802_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [9:0] SBMux_C24_N23804_O_3_C_7_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C24_N23804_O_3_C_7_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C24_N23804_O_3_C_7_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C24_N23804_O_3_C_7_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C24_N23804_O_3_C_7_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C24_N23804_O_3_C_7_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C24_N23804_O_3_C_7_io_arst; // @[TileFull.scala 141:27]
  wire [7:0] SBMux_C32_N23806_O_3_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C32_N23806_O_3_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C32_N23806_O_3_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C32_N23806_O_3_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C32_N23806_O_3_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C32_N23806_O_3_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C32_N23806_O_3_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [7:0] SBMux_C40_N23808_O_3_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C40_N23808_O_3_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C40_N23808_O_3_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C40_N23808_O_3_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C40_N23808_O_3_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C40_N23808_O_3_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C40_N23808_O_3_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C48_N23810_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C48_N23810_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C48_N23810_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C48_N23810_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C48_N23810_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C48_N23810_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C48_N23810_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C56_N23812_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C56_N23812_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C56_N23812_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C56_N23812_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C56_N23812_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C56_N23812_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C56_N23812_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C64_N23814_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C64_N23814_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C64_N23814_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C64_N23814_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C64_N23814_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C64_N23814_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C64_N23814_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [9:0] SBMux_C72_N23816_O_3_C_7_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C72_N23816_O_3_C_7_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C72_N23816_O_3_C_7_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C72_N23816_O_3_C_7_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C72_N23816_O_3_C_7_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C72_N23816_O_3_C_7_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C72_N23816_O_3_C_7_io_arst; // @[TileFull.scala 141:27]
  wire [7:0] SBMux_C80_N23818_O_2_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C80_N23818_O_2_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C80_N23818_O_2_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C80_N23818_O_2_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C80_N23818_O_2_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C80_N23818_O_2_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C80_N23818_O_2_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [7:0] SBMux_C88_N23820_O_3_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C88_N23820_O_3_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C88_N23820_O_3_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C88_N23820_O_3_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C88_N23820_O_3_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C88_N23820_O_3_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C88_N23820_O_3_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [6:0] SBMux_C96_N23822_O_2_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C96_N23822_O_2_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C96_N23822_O_2_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C96_N23822_O_2_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C96_N23822_O_2_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C96_N23822_O_2_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C96_N23822_O_2_C_5_io_arst; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N23824_O_0_C_1_io_in; // @[TileFull.scala 141:27]
  wire [1:0] SBMux_C100_N23824_O_0_C_1_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N23824_O_0_C_1_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N23824_O_0_C_1_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N23824_O_0_C_1_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N23824_O_0_C_1_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N23824_O_0_C_1_io_arst; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N23826_O_0_C_1_io_in; // @[TileFull.scala 141:27]
  wire [1:0] SBMux_C104_N23826_O_0_C_1_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N23826_O_0_C_1_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N23826_O_0_C_1_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N23826_O_0_C_1_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N23826_O_0_C_1_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N23826_O_0_C_1_io_arst; // @[TileFull.scala 141:27]
  wire [9:0] SBMux_C1_N30079_O_4_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C1_N30079_O_4_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C1_N30079_O_4_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C1_N30079_O_4_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C1_N30079_O_4_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C1_N30079_O_4_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C1_N30079_O_4_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [10:0] SBMux_C9_N30087_O_4_C_7_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C9_N30087_O_4_C_7_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C9_N30087_O_4_C_7_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C9_N30087_O_4_C_7_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C9_N30087_O_4_C_7_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C9_N30087_O_4_C_7_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C9_N30087_O_4_C_7_io_arst; // @[TileFull.scala 141:27]
  wire [9:0] SBMux_C17_N30095_O_3_C_7_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C17_N30095_O_3_C_7_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C17_N30095_O_3_C_7_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C17_N30095_O_3_C_7_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C17_N30095_O_3_C_7_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C17_N30095_O_3_C_7_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C17_N30095_O_3_C_7_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C25_N30103_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C25_N30103_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C25_N30103_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C25_N30103_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C25_N30103_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C25_N30103_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C25_N30103_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [6:0] SBMux_C33_N30111_O_3_C_4_io_in; // @[TileFull.scala 141:27]
  wire [2:0] SBMux_C33_N30111_O_3_C_4_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C33_N30111_O_3_C_4_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C33_N30111_O_3_C_4_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C33_N30111_O_3_C_4_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C33_N30111_O_3_C_4_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C33_N30111_O_3_C_4_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C41_N30119_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C41_N30119_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C41_N30119_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C41_N30119_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C41_N30119_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C41_N30119_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C41_N30119_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C49_N30127_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C49_N30127_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C49_N30127_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C49_N30127_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C49_N30127_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C49_N30127_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C49_N30127_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C57_N30135_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C57_N30135_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C57_N30135_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C57_N30135_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C57_N30135_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C57_N30135_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C57_N30135_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C65_N30143_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C65_N30143_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C65_N30143_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C65_N30143_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C65_N30143_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C65_N30143_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C65_N30143_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C73_N30151_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C73_N30151_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C73_N30151_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C73_N30151_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C73_N30151_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C73_N30151_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C73_N30151_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C81_N30159_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C81_N30159_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C81_N30159_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C81_N30159_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C81_N30159_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C81_N30159_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C81_N30159_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C89_N30167_O_4_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C89_N30167_O_4_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C89_N30167_O_4_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C89_N30167_O_4_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C89_N30167_O_4_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C89_N30167_O_4_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C89_N30167_O_4_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C97_N30175_O_4_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C97_N30175_O_4_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C97_N30175_O_4_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C97_N30175_O_4_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C97_N30175_O_4_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C97_N30175_O_4_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C97_N30175_O_4_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [4:0] SBMux_C101_N30179_O_4_C_1_io_in; // @[TileFull.scala 141:27]
  wire [2:0] SBMux_C101_N30179_O_4_C_1_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N30179_O_4_C_1_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N30179_O_4_C_1_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N30179_O_4_C_1_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N30179_O_4_C_1_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C101_N30179_O_4_C_1_io_arst; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C105_N30183_O_3_C_1_io_in; // @[TileFull.scala 141:27]
  wire [2:0] SBMux_C105_N30183_O_3_C_1_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N30183_O_3_C_1_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N30183_O_3_C_1_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N30183_O_3_C_1_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N30183_O_3_C_1_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C105_N30183_O_3_C_1_io_arst; // @[TileFull.scala 141:27]
  wire [9:0] SBMux_C0_N30186_O_4_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C0_N30186_O_4_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C0_N30186_O_4_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C0_N30186_O_4_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C0_N30186_O_4_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C0_N30186_O_4_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C0_N30186_O_4_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C8_N30188_O_4_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C8_N30188_O_4_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C8_N30188_O_4_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C8_N30188_O_4_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C8_N30188_O_4_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C8_N30188_O_4_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C8_N30188_O_4_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [9:0] SBMux_C16_N30190_O_3_C_7_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C16_N30190_O_3_C_7_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C16_N30190_O_3_C_7_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C16_N30190_O_3_C_7_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C16_N30190_O_3_C_7_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C16_N30190_O_3_C_7_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C16_N30190_O_3_C_7_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C24_N30192_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C24_N30192_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C24_N30192_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C24_N30192_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C24_N30192_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C24_N30192_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C24_N30192_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C32_N30194_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C32_N30194_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C32_N30194_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C32_N30194_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C32_N30194_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C32_N30194_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C32_N30194_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [7:0] SBMux_C40_N30196_O_3_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C40_N30196_O_3_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C40_N30196_O_3_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C40_N30196_O_3_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C40_N30196_O_3_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C40_N30196_O_3_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C40_N30196_O_3_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C48_N30198_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C48_N30198_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C48_N30198_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C48_N30198_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C48_N30198_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C48_N30198_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C48_N30198_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C56_N30200_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C56_N30200_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C56_N30200_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C56_N30200_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C56_N30200_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C56_N30200_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C56_N30200_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [9:0] SBMux_C64_N30202_O_3_C_7_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C64_N30202_O_3_C_7_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C64_N30202_O_3_C_7_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C64_N30202_O_3_C_7_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C64_N30202_O_3_C_7_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C64_N30202_O_3_C_7_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C64_N30202_O_3_C_7_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C72_N30204_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C72_N30204_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C72_N30204_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C72_N30204_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C72_N30204_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C72_N30204_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C72_N30204_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C80_N30206_O_3_C_6_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C80_N30206_O_3_C_6_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C80_N30206_O_3_C_6_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C80_N30206_O_3_C_6_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C80_N30206_O_3_C_6_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C80_N30206_O_3_C_6_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C80_N30206_O_3_C_6_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C88_N30208_O_4_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C88_N30208_O_4_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C88_N30208_O_4_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C88_N30208_O_4_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C88_N30208_O_4_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C88_N30208_O_4_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C88_N30208_O_4_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [8:0] SBMux_C96_N30210_O_4_C_5_io_in; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C96_N30210_O_4_C_5_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C96_N30210_O_4_C_5_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C96_N30210_O_4_C_5_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C96_N30210_O_4_C_5_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C96_N30210_O_4_C_5_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C96_N30210_O_4_C_5_io_arst; // @[TileFull.scala 141:27]
  wire [4:0] SBMux_C100_N30212_O_4_C_1_io_in; // @[TileFull.scala 141:27]
  wire [2:0] SBMux_C100_N30212_O_4_C_1_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N30212_O_4_C_1_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N30212_O_4_C_1_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N30212_O_4_C_1_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N30212_O_4_C_1_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C100_N30212_O_4_C_1_io_arst; // @[TileFull.scala 141:27]
  wire [3:0] SBMux_C104_N30214_O_3_C_1_io_in; // @[TileFull.scala 141:27]
  wire [2:0] SBMux_C104_N30214_O_3_C_1_io_config; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N30214_O_3_C_1_io_out; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N30214_O_3_C_1_io_loopBreak; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N30214_O_3_C_1_io_ioGndBle; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N30214_O_3_C_1_io_cnstClk; // @[TileFull.scala 141:27]
  wire  SBMux_C104_N30214_O_3_C_1_io_arst; // @[TileFull.scala 141:27]
  wire  _CBMux_IPIN0_N14762_io_in_WIRE_1 = SBMux_C1_N30079_O_4_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN0_N14762_io_in_WIRE_5 = SBMux_C9_N30087_O_4_C_7_io_out; // @[TileFull.scala 170:{37,37}]
  wire [6:0] CBMux_IPIN0_N14762_io_in_lo_lo = {IN_CHANY_N30094_16,_CBMux_IPIN0_N14762_io_in_WIRE_5,IN_CHANY_N30086_8,
    IN_CHANY_N30081_3,IN_CHANY_N30080_2,_CBMux_IPIN0_N14762_io_in_WIRE_1,IN_CHANY_N30078_0}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN0_N14762_io_in_WIRE_9 = SBMux_C25_N30103_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN0_N14762_io_in_WIRE_7 = SBMux_C17_N30095_O_3_C_7_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN0_N14762_io_in_WIRE_11 = SBMux_C33_N30111_O_3_C_4_io_out; // @[TileFull.scala 170:{37,37}]
  wire [13:0] CBMux_IPIN0_N14762_io_in_lo = {IN_CHANY_N30125_47,IN_CHANY_N30124_46,_CBMux_IPIN0_N14762_io_in_WIRE_11,
    IN_CHANY_N30110_32,_CBMux_IPIN0_N14762_io_in_WIRE_9,IN_CHANY_N30102_24,_CBMux_IPIN0_N14762_io_in_WIRE_7,
    CBMux_IPIN0_N14762_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN0_N14762_io_in_hi_lo = {IN_CHANY_N30156_78,IN_CHANY_N30149_71,IN_CHANY_N30148_70,
    IN_CHANY_N30141_63,IN_CHANY_N30140_62,IN_CHANY_N30133_55,IN_CHANY_N30132_54}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN0_N14762_io_in_hi = {IN_CHANY_N30181_103,IN_CHANY_N30180_102,IN_CHANY_N30173_95,
    IN_CHANY_N30172_94,IN_CHANY_N30165_87,IN_CHANY_N30164_86,IN_CHANY_N30157_79,CBMux_IPIN0_N14762_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN1_N14763_io_in_lo_lo = {IN_CHANY_N30104_26,IN_CHANY_N30097_19,IN_CHANY_N30096_18,
    IN_CHANY_N30089_11,IN_CHANY_N30088_10,IN_CHANY_N30083_5,IN_CHANY_N30082_4}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN1_N14763_io_in_WIRE_11 = SBMux_C41_N30119_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire [13:0] CBMux_IPIN1_N14763_io_in_lo = {IN_CHANY_N30121_43,IN_CHANY_N30120_42,_CBMux_IPIN1_N14763_io_in_WIRE_11,
    IN_CHANY_N30118_40,IN_CHANY_N30113_35,IN_CHANY_N30112_34,IN_CHANY_N30105_27,CBMux_IPIN1_N14763_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN1_N14763_io_in_WIRE_15 = SBMux_C49_N30127_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN1_N14763_io_in_WIRE_17 = SBMux_C57_N30135_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN1_N14763_io_in_WIRE_19 = SBMux_C65_N30143_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire [6:0] CBMux_IPIN1_N14763_io_in_hi_lo = {IN_CHANY_N30150_72,_CBMux_IPIN1_N14763_io_in_WIRE_19,IN_CHANY_N30142_64,
    _CBMux_IPIN1_N14763_io_in_WIRE_17,IN_CHANY_N30134_56,_CBMux_IPIN1_N14763_io_in_WIRE_15,IN_CHANY_N30126_48}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN1_N14763_io_in_WIRE_23 = SBMux_C89_N30167_O_4_C_5_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN1_N14763_io_in_WIRE_21 = SBMux_C73_N30151_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN1_N14763_io_in_WIRE_25 = SBMux_C97_N30175_O_4_C_5_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN1_N14763_io_in_WIRE_27 = SBMux_C101_N30179_O_4_C_1_io_out; // @[TileFull.scala 170:{37,37}]
  wire [13:0] CBMux_IPIN1_N14763_io_in_hi = {_CBMux_IPIN1_N14763_io_in_WIRE_27,IN_CHANY_N30178_100,
    _CBMux_IPIN1_N14763_io_in_WIRE_25,IN_CHANY_N30174_96,_CBMux_IPIN1_N14763_io_in_WIRE_23,IN_CHANY_N30166_88,
    _CBMux_IPIN1_N14763_io_in_WIRE_21,CBMux_IPIN1_N14763_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN2_N14764_io_in_lo_lo = {IN_CHANY_N30106_28,IN_CHANY_N30099_21,IN_CHANY_N30098_20,
    IN_CHANY_N30091_13,IN_CHANY_N30090_12,IN_CHANY_N30085_7,IN_CHANY_N30084_6}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN2_N14764_io_in_lo = {IN_CHANY_N30129_51,IN_CHANY_N30128_50,IN_CHANY_N30123_45,IN_CHANY_N30122_44
    ,IN_CHANY_N30115_37,IN_CHANY_N30114_36,IN_CHANY_N30107_29,CBMux_IPIN2_N14764_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN2_N14764_io_in_hi_lo = {IN_CHANY_N30160_82,IN_CHANY_N30153_75,IN_CHANY_N30152_74,
    IN_CHANY_N30145_67,IN_CHANY_N30144_66,IN_CHANY_N30137_59,IN_CHANY_N30136_58}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN2_N14764_io_in_hi = {IN_CHANY_N30185_107,IN_CHANY_N30184_106,IN_CHANY_N30177_99,
    IN_CHANY_N30176_98,IN_CHANY_N30169_91,IN_CHANY_N30168_90,IN_CHANY_N30161_83,CBMux_IPIN2_N14764_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN3_N14765_io_in_lo_lo = {IN_CHANY_N30108_30,IN_CHANY_N30101_23,IN_CHANY_N30100_22,
    IN_CHANY_N30093_15,IN_CHANY_N30092_14,IN_CHANY_N30085_7,IN_CHANY_N30084_6}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN3_N14765_io_in_lo = {IN_CHANY_N30131_53,IN_CHANY_N30130_52,IN_CHANY_N30125_47,IN_CHANY_N30124_46
    ,IN_CHANY_N30117_39,IN_CHANY_N30116_38,IN_CHANY_N30109_31,CBMux_IPIN3_N14765_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN3_N14765_io_in_hi_lo = {IN_CHANY_N30158_80,IN_CHANY_N30155_77,IN_CHANY_N30154_76,
    IN_CHANY_N30147_69,IN_CHANY_N30146_68,IN_CHANY_N30139_61,IN_CHANY_N30138_60}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN3_N14765_io_in_WIRE_21 = SBMux_C81_N30159_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN3_N14765_io_in_WIRE_27 = SBMux_C105_N30183_O_3_C_1_io_out; // @[TileFull.scala 170:{37,37}]
  wire [13:0] CBMux_IPIN3_N14765_io_in_hi = {_CBMux_IPIN3_N14765_io_in_WIRE_27,IN_CHANY_N30182_104,IN_CHANY_N30171_93,
    IN_CHANY_N30170_92,IN_CHANY_N30163_85,IN_CHANY_N30162_84,_CBMux_IPIN3_N14765_io_in_WIRE_21,
    CBMux_IPIN3_N14765_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN4_N14766_io_in_lo = {_CBMux_IPIN1_N14763_io_in_WIRE_11,IN_CHANY_N30118_40,
    _CBMux_IPIN0_N14762_io_in_WIRE_11,IN_CHANY_N30110_32,_CBMux_IPIN0_N14762_io_in_WIRE_9,IN_CHANY_N30102_24,
    _CBMux_IPIN0_N14762_io_in_WIRE_7,CBMux_IPIN0_N14762_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN4_N14766_io_in_hi = {_CBMux_IPIN3_N14765_io_in_WIRE_27,IN_CHANY_N30182_104,IN_CHANY_N30171_93,
    IN_CHANY_N30170_92,IN_CHANY_N30163_85,IN_CHANY_N30162_84,IN_CHANY_N30157_79,CBMux_IPIN0_N14762_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN5_N14767_io_in_lo = {_CBMux_IPIN1_N14763_io_in_WIRE_15,IN_CHANY_N30126_48,IN_CHANY_N30121_43,
    IN_CHANY_N30120_42,IN_CHANY_N30113_35,IN_CHANY_N30112_34,IN_CHANY_N30105_27,CBMux_IPIN1_N14763_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN5_N14767_io_in_hi_lo = {IN_CHANY_N30150_72,_CBMux_IPIN1_N14763_io_in_WIRE_19,IN_CHANY_N30142_64,
    _CBMux_IPIN1_N14763_io_in_WIRE_17,IN_CHANY_N30134_56,IN_CHANY_N30129_51,IN_CHANY_N30128_50}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN5_N14767_io_in_hi = {IN_CHANY_N30181_103,IN_CHANY_N30180_102,IN_CHANY_N30173_95,
    IN_CHANY_N30172_94,IN_CHANY_N30165_87,IN_CHANY_N30164_86,_CBMux_IPIN1_N14763_io_in_WIRE_21,
    CBMux_IPIN5_N14767_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN6_N14768_io_in_lo = {IN_CHANY_N30131_53,IN_CHANY_N30130_52,IN_CHANY_N30123_45,IN_CHANY_N30122_44
    ,IN_CHANY_N30115_37,IN_CHANY_N30114_36,IN_CHANY_N30107_29,CBMux_IPIN2_N14764_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN6_N14768_io_in_hi = {_CBMux_IPIN1_N14763_io_in_WIRE_27,IN_CHANY_N30178_100,
    _CBMux_IPIN1_N14763_io_in_WIRE_25,IN_CHANY_N30174_96,_CBMux_IPIN1_N14763_io_in_WIRE_23,IN_CHANY_N30166_88,
    IN_CHANY_N30161_83,CBMux_IPIN2_N14764_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN7_N14769_io_in_lo = {IN_CHANY_N30131_53,IN_CHANY_N30130_52,IN_CHANY_N30123_45,IN_CHANY_N30122_44
    ,IN_CHANY_N30117_39,IN_CHANY_N30116_38,IN_CHANY_N30109_31,CBMux_IPIN3_N14765_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN7_N14769_io_in_hi = {IN_CHANY_N30185_107,IN_CHANY_N30184_106,IN_CHANY_N30177_99,
    IN_CHANY_N30176_98,IN_CHANY_N30169_91,IN_CHANY_N30168_90,_CBMux_IPIN3_N14765_io_in_WIRE_21,
    CBMux_IPIN3_N14765_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN8_N14770_io_in_lo_lo = {IN_CHANY_N30108_30,IN_CHANY_N30101_23,IN_CHANY_N30100_22,
    _CBMux_IPIN0_N14762_io_in_WIRE_5,IN_CHANY_N30086_8,_CBMux_IPIN0_N14762_io_in_WIRE_1,IN_CHANY_N30078_0}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN8_N14770_io_in_lo = {IN_CHANY_N30133_55,IN_CHANY_N30132_54,IN_CHANY_N30125_47,IN_CHANY_N30124_46
    ,IN_CHANY_N30117_39,IN_CHANY_N30116_38,IN_CHANY_N30109_31,CBMux_IPIN8_N14770_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN9_N14771_io_in_lo_lo = {IN_CHANY_N30096_18,_CBMux_IPIN0_N14762_io_in_WIRE_7,IN_CHANY_N30094_16,
    IN_CHANY_N30089_11,IN_CHANY_N30088_10,IN_CHANY_N30081_3,IN_CHANY_N30080_2}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN9_N14771_io_in_lo = {_CBMux_IPIN1_N14763_io_in_WIRE_11,IN_CHANY_N30118_40,
    _CBMux_IPIN0_N14762_io_in_WIRE_11,IN_CHANY_N30110_32,_CBMux_IPIN0_N14762_io_in_WIRE_9,IN_CHANY_N30102_24,
    IN_CHANY_N30097_19,CBMux_IPIN9_N14771_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN9_N14771_io_in_hi_lo = {IN_CHANY_N30156_78,IN_CHANY_N30149_71,IN_CHANY_N30148_70,
    IN_CHANY_N30141_63,IN_CHANY_N30140_62,_CBMux_IPIN1_N14763_io_in_WIRE_15,IN_CHANY_N30126_48}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN9_N14771_io_in_hi = {_CBMux_IPIN3_N14765_io_in_WIRE_27,IN_CHANY_N30182_104,IN_CHANY_N30171_93,
    IN_CHANY_N30170_92,IN_CHANY_N30163_85,IN_CHANY_N30162_84,IN_CHANY_N30157_79,CBMux_IPIN9_N14771_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN10_N14772_io_in_lo_lo = {IN_CHANY_N30104_26,IN_CHANY_N30099_21,IN_CHANY_N30098_20,
    IN_CHANY_N30091_13,IN_CHANY_N30090_12,IN_CHANY_N30083_5,IN_CHANY_N30082_4}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN10_N14772_io_in_lo = {IN_CHANY_N30129_51,IN_CHANY_N30128_50,IN_CHANY_N30121_43,
    IN_CHANY_N30120_42,IN_CHANY_N30113_35,IN_CHANY_N30112_34,IN_CHANY_N30105_27,CBMux_IPIN10_N14772_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN10_N14772_io_in_hi_lo = {IN_CHANY_N30150_72,_CBMux_IPIN1_N14763_io_in_WIRE_19,IN_CHANY_N30142_64,
    IN_CHANY_N30137_59,IN_CHANY_N30136_58,_CBMux_IPIN1_N14763_io_in_WIRE_17,IN_CHANY_N30134_56}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN10_N14772_io_in_hi = {IN_CHANY_N30181_103,IN_CHANY_N30180_102,IN_CHANY_N30173_95,
    IN_CHANY_N30172_94,IN_CHANY_N30165_87,IN_CHANY_N30164_86,_CBMux_IPIN1_N14763_io_in_WIRE_21,
    CBMux_IPIN10_N14772_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN11_N14773_io_in_lo_lo = {IN_CHANY_N30106_28,IN_CHANY_N30099_21,IN_CHANY_N30098_20,
    IN_CHANY_N30093_15,IN_CHANY_N30092_14,IN_CHANY_N30085_7,IN_CHANY_N30084_6}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN11_N14773_io_in_lo = {IN_CHANY_N30131_53,IN_CHANY_N30130_52,IN_CHANY_N30123_45,
    IN_CHANY_N30122_44,IN_CHANY_N30115_37,IN_CHANY_N30114_36,IN_CHANY_N30107_29,CBMux_IPIN11_N14773_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN12_N14774_io_in_lo_lo = {IN_CHANY_N30108_30,IN_CHANY_N30101_23,IN_CHANY_N30100_22,
    IN_CHANY_N30093_15,IN_CHANY_N30092_14,_CBMux_IPIN0_N14762_io_in_WIRE_1,IN_CHANY_N30078_0}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN12_N14774_io_in_lo = {IN_CHANY_N30133_55,IN_CHANY_N30132_54,IN_CHANY_N30125_47,
    IN_CHANY_N30124_46,IN_CHANY_N30117_39,IN_CHANY_N30116_38,IN_CHANY_N30109_31,CBMux_IPIN12_N14774_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN12_N14774_io_in_hi = {_CBMux_IPIN1_N14763_io_in_WIRE_27,IN_CHANY_N30178_100,
    _CBMux_IPIN1_N14763_io_in_WIRE_25,IN_CHANY_N30174_96,_CBMux_IPIN1_N14763_io_in_WIRE_23,IN_CHANY_N30166_88,
    _CBMux_IPIN3_N14765_io_in_WIRE_21,CBMux_IPIN3_N14765_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN13_N14775_io_in_lo_lo = {IN_CHANY_N30094_16,IN_CHANY_N30089_11,IN_CHANY_N30088_10,
    _CBMux_IPIN0_N14762_io_in_WIRE_5,IN_CHANY_N30086_8,IN_CHANY_N30081_3,IN_CHANY_N30080_2}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN13_N14775_io_in_lo = {_CBMux_IPIN1_N14763_io_in_WIRE_11,IN_CHANY_N30118_40,
    _CBMux_IPIN0_N14762_io_in_WIRE_11,IN_CHANY_N30110_32,_CBMux_IPIN0_N14762_io_in_WIRE_9,IN_CHANY_N30102_24,
    _CBMux_IPIN0_N14762_io_in_WIRE_7,CBMux_IPIN13_N14775_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN13_N14775_io_in_hi = {IN_CHANY_N30185_107,IN_CHANY_N30184_106,IN_CHANY_N30177_99,
    IN_CHANY_N30176_98,IN_CHANY_N30169_91,IN_CHANY_N30168_90,IN_CHANY_N30157_79,CBMux_IPIN9_N14771_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN14_N14776_io_in_lo_lo = {IN_CHANY_N30104_26,IN_CHANY_N30097_19,IN_CHANY_N30096_18,
    IN_CHANY_N30091_13,IN_CHANY_N30090_12,IN_CHANY_N30083_5,IN_CHANY_N30082_4}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN14_N14776_io_in_lo = {_CBMux_IPIN1_N14763_io_in_WIRE_15,IN_CHANY_N30126_48,IN_CHANY_N30121_43,
    IN_CHANY_N30120_42,IN_CHANY_N30113_35,IN_CHANY_N30112_34,IN_CHANY_N30105_27,CBMux_IPIN14_N14776_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN14_N14776_io_in_hi = {_CBMux_IPIN3_N14765_io_in_WIRE_27,IN_CHANY_N30182_104,IN_CHANY_N30171_93,
    IN_CHANY_N30170_92,IN_CHANY_N30163_85,IN_CHANY_N30162_84,_CBMux_IPIN1_N14763_io_in_WIRE_21,
    CBMux_IPIN5_N14767_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN15_N14777_io_in_lo_lo = {IN_CHANY_N30106_28,IN_CHANY_N30099_21,IN_CHANY_N30098_20,
    IN_CHANY_N30091_13,IN_CHANY_N30090_12,IN_CHANY_N30083_5,IN_CHANY_N30082_4}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN15_N14777_io_in_lo = {IN_CHANY_N30129_51,IN_CHANY_N30128_50,IN_CHANY_N30121_43,
    IN_CHANY_N30120_42,IN_CHANY_N30115_37,IN_CHANY_N30114_36,IN_CHANY_N30107_29,CBMux_IPIN15_N14777_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN15_N14777_io_in_hi = {IN_CHANY_N30181_103,IN_CHANY_N30180_102,IN_CHANY_N30173_95,
    IN_CHANY_N30172_94,IN_CHANY_N30165_87,IN_CHANY_N30164_86,IN_CHANY_N30161_83,CBMux_IPIN2_N14764_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN16_N14778_io_in_WIRE_1 = SBMux_C1_N23683_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN16_N14778_io_in_WIRE_3 = SBMux_C9_N23685_O_3_C_7_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN16_N14778_io_in_WIRE_5 = SBMux_C17_N23687_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire [6:0] CBMux_IPIN16_N14778_io_in_lo_lo = {IN_CHANX_N23688_24,_CBMux_IPIN16_N14778_io_in_WIRE_5,IN_CHANX_N23686_16,
    _CBMux_IPIN16_N14778_io_in_WIRE_3,IN_CHANX_N23684_8,_CBMux_IPIN16_N14778_io_in_WIRE_1,IN_CHANX_N23682_0}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN16_N14778_io_in_WIRE_9 = SBMux_C33_N23691_O_3_C_7_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN16_N14778_io_in_WIRE_7 = SBMux_C25_N23689_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire [13:0] CBMux_IPIN16_N14778_io_in_lo = {IN_CHANX_N23781_47,IN_CHANX_N23780_46,IN_CHANX_N23713_3,IN_CHANX_N23712_2,
    _CBMux_IPIN16_N14778_io_in_WIRE_9,IN_CHANX_N23690_32,_CBMux_IPIN16_N14778_io_in_WIRE_7,
    CBMux_IPIN16_N14778_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN16_N14778_io_in_hi_lo = {IN_CHANX_N23788_78,IN_CHANX_N23787_71,IN_CHANX_N23786_70,
    IN_CHANX_N23785_63,IN_CHANX_N23784_62,IN_CHANX_N23783_55,IN_CHANX_N23782_54}; // @[TileFull.scala 175:8]
  wire [13:0] CBMux_IPIN16_N14778_io_in_hi = {IN_CHANX_N23795_103,IN_CHANX_N23794_102,IN_CHANX_N23793_95,
    IN_CHANX_N23792_94,IN_CHANX_N23791_87,IN_CHANX_N23790_86,IN_CHANX_N23789_79,CBMux_IPIN16_N14778_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN17_N14779_io_in_WIRE_1 = SBMux_C41_N23693_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN17_N14779_io_in_WIRE_3 = SBMux_C49_N23695_O_3_C_5_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN17_N14779_io_in_WIRE_5 = SBMux_C57_N23697_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire [6:0] CBMux_IPIN17_N14779_io_in_lo_lo = {IN_CHANX_N23698_64,_CBMux_IPIN17_N14779_io_in_WIRE_5,IN_CHANX_N23696_56,
    _CBMux_IPIN17_N14779_io_in_WIRE_3,IN_CHANX_N23694_48,_CBMux_IPIN17_N14779_io_in_WIRE_1,IN_CHANX_N23692_40}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN17_N14779_io_in_WIRE_9 = SBMux_C73_N23701_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN17_N14779_io_in_WIRE_7 = SBMux_C65_N23699_O_3_C_6_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN17_N14779_io_in_WIRE_11 = SBMux_C89_N23705_O_3_C_5_io_out; // @[TileFull.scala 170:{37,37}]
  wire  _CBMux_IPIN17_N14779_io_in_WIRE_13 = SBMux_C97_N23707_O_2_C_5_io_out; // @[TileFull.scala 170:{37,37}]
  wire [13:0] CBMux_IPIN17_N14779_io_in_lo = {_CBMux_IPIN17_N14779_io_in_WIRE_13,IN_CHANX_N23706_96,
    _CBMux_IPIN17_N14779_io_in_WIRE_11,IN_CHANX_N23704_88,_CBMux_IPIN17_N14779_io_in_WIRE_9,IN_CHANX_N23700_72,
    _CBMux_IPIN17_N14779_io_in_WIRE_7,CBMux_IPIN17_N14779_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [6:0] CBMux_IPIN17_N14779_io_in_hi_lo = {IN_CHANX_N23720_34,IN_CHANX_N23719_27,IN_CHANX_N23718_26,
    IN_CHANX_N23717_19,IN_CHANX_N23716_18,IN_CHANX_N23715_11,IN_CHANX_N23714_10}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN17_N14779_io_in_WIRE_27 = SBMux_C101_N23767_O_0_C_1_io_out; // @[TileFull.scala 170:{37,37}]
  wire [13:0] CBMux_IPIN17_N14779_io_in_hi = {_CBMux_IPIN17_N14779_io_in_WIRE_27,IN_CHANX_N23766_100,IN_CHANX_N23743_5,
    IN_CHANX_N23742_4,IN_CHANX_N23723_43,IN_CHANX_N23722_42,IN_CHANX_N23721_35,CBMux_IPIN17_N14779_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN18_N14780_io_in_lo_lo = {IN_CHANX_N23729_67,IN_CHANX_N23728_66,IN_CHANX_N23727_59,
    IN_CHANX_N23726_58,IN_CHANX_N23725_51,IN_CHANX_N23724_50}; // @[TileFull.scala 175:8]
  wire [11:0] CBMux_IPIN18_N14780_io_in_lo = {IN_CHANX_N23745_13,IN_CHANX_N23744_12,IN_CHANX_N23733_83,
    IN_CHANX_N23732_82,IN_CHANX_N23731_75,IN_CHANX_N23730_74,CBMux_IPIN18_N14780_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN18_N14780_io_in_hi_lo = {IN_CHANX_N23751_37,IN_CHANX_N23750_36,IN_CHANX_N23749_29,
    IN_CHANX_N23748_28,IN_CHANX_N23747_21,IN_CHANX_N23746_20}; // @[TileFull.scala 175:8]
  wire [11:0] CBMux_IPIN18_N14780_io_in_hi = {IN_CHANX_N23797_107,IN_CHANX_N23796_106,IN_CHANX_N23771_7,
    IN_CHANX_N23770_6,IN_CHANX_N23753_45,IN_CHANX_N23752_44,CBMux_IPIN18_N14780_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN19_N14781_io_in_WIRE_1 = SBMux_C81_N23703_O_2_C_5_io_out; // @[TileFull.scala 170:{37,37}]
  wire [5:0] CBMux_IPIN19_N14781_io_in_lo_lo = {IN_CHANX_N23755_53,IN_CHANX_N23754_52,IN_CHANX_N23753_45,
    IN_CHANX_N23752_44,_CBMux_IPIN19_N14781_io_in_WIRE_1,IN_CHANX_N23702_80}; // @[TileFull.scala 175:8]
  wire [11:0] CBMux_IPIN19_N14781_io_in_lo = {IN_CHANX_N23761_77,IN_CHANX_N23760_76,IN_CHANX_N23759_69,
    IN_CHANX_N23758_68,IN_CHANX_N23757_61,IN_CHANX_N23756_60,CBMux_IPIN19_N14781_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire  _CBMux_IPIN19_N14781_io_in_WIRE_13 = SBMux_C105_N23769_O_0_C_1_io_out; // @[TileFull.scala 170:{37,37}]
  wire [5:0] CBMux_IPIN19_N14781_io_in_hi_lo = {IN_CHANX_N23773_15,IN_CHANX_N23772_14,IN_CHANX_N23771_7,
    IN_CHANX_N23770_6,_CBMux_IPIN19_N14781_io_in_WIRE_13,IN_CHANX_N23768_104}; // @[TileFull.scala 175:8]
  wire [11:0] CBMux_IPIN19_N14781_io_in_hi = {IN_CHANX_N23779_39,IN_CHANX_N23778_38,IN_CHANX_N23777_31,
    IN_CHANX_N23776_30,IN_CHANX_N23775_23,IN_CHANX_N23774_22,CBMux_IPIN19_N14781_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN20_N14782_io_in_lo_lo = {IN_CHANX_N23754_52,_CBMux_IPIN19_N14781_io_in_WIRE_1,IN_CHANX_N23702_80,
    _CBMux_IPIN16_N14778_io_in_WIRE_1,IN_CHANX_N23682_0}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN20_N14782_io_in_lo = {IN_CHANX_N23760_76,IN_CHANX_N23759_69,IN_CHANX_N23758_68,
    IN_CHANX_N23757_61,IN_CHANX_N23756_60,IN_CHANX_N23755_53,CBMux_IPIN20_N14782_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN20_N14782_io_in_hi_lo = {IN_CHANX_N23775_23,IN_CHANX_N23774_22,IN_CHANX_N23773_15,
    IN_CHANX_N23772_14,IN_CHANX_N23761_77}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN20_N14782_io_in_hi = {IN_CHANX_N23781_47,IN_CHANX_N23780_46,IN_CHANX_N23779_39,
    IN_CHANX_N23778_38,IN_CHANX_N23777_31,IN_CHANX_N23776_30,CBMux_IPIN20_N14782_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN21_N14783_io_in_lo_lo = {_CBMux_IPIN16_N14778_io_in_WIRE_7,IN_CHANX_N23688_24,
    _CBMux_IPIN16_N14778_io_in_WIRE_5,IN_CHANX_N23686_16,_CBMux_IPIN16_N14778_io_in_WIRE_3,IN_CHANX_N23684_8}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN21_N14783_io_in_lo = {IN_CHANX_N23714_10,IN_CHANX_N23713_3,IN_CHANX_N23712_2,
    _CBMux_IPIN17_N14779_io_in_WIRE_1,IN_CHANX_N23692_40,_CBMux_IPIN16_N14778_io_in_WIRE_9,IN_CHANX_N23690_32,
    CBMux_IPIN21_N14783_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN21_N14783_io_in_hi_lo = {IN_CHANX_N23786_70,IN_CHANX_N23785_63,IN_CHANX_N23784_62,
    IN_CHANX_N23783_55,IN_CHANX_N23782_54,IN_CHANX_N23715_11}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN21_N14783_io_in_hi = {IN_CHANX_N23793_95,IN_CHANX_N23792_94,IN_CHANX_N23791_87,
    IN_CHANX_N23790_86,IN_CHANX_N23789_79,IN_CHANX_N23788_78,IN_CHANX_N23787_71,CBMux_IPIN21_N14783_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN22_N14784_io_in_lo_lo = {_CBMux_IPIN17_N14779_io_in_WIRE_7,IN_CHANX_N23698_64,
    _CBMux_IPIN17_N14779_io_in_WIRE_5,IN_CHANX_N23696_56,_CBMux_IPIN17_N14779_io_in_WIRE_3,IN_CHANX_N23694_48}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN22_N14784_io_in_lo = {IN_CHANX_N23716_18,_CBMux_IPIN17_N14779_io_in_WIRE_13,IN_CHANX_N23706_96,
    _CBMux_IPIN17_N14779_io_in_WIRE_11,IN_CHANX_N23704_88,_CBMux_IPIN17_N14779_io_in_WIRE_9,IN_CHANX_N23700_72,
    CBMux_IPIN22_N14784_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN22_N14784_io_in_hi_lo = {IN_CHANX_N23722_42,IN_CHANX_N23721_35,IN_CHANX_N23720_34,
    IN_CHANX_N23719_27,IN_CHANX_N23718_26,IN_CHANX_N23717_19}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN22_N14784_io_in_hi = {IN_CHANX_N23745_13,IN_CHANX_N23744_12,IN_CHANX_N23743_5,IN_CHANX_N23742_4,
    IN_CHANX_N23725_51,IN_CHANX_N23724_50,IN_CHANX_N23723_43,CBMux_IPIN22_N14784_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN23_N14785_io_in_lo_lo = {IN_CHANX_N23730_74,IN_CHANX_N23729_67,IN_CHANX_N23728_66,
    IN_CHANX_N23727_59,IN_CHANX_N23726_58}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN23_N14785_io_in_lo = {IN_CHANX_N23746_20,IN_CHANX_N23745_13,IN_CHANX_N23744_12,
    IN_CHANX_N23733_83,IN_CHANX_N23732_82,IN_CHANX_N23731_75,CBMux_IPIN23_N14785_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN23_N14785_io_in_hi_lo = {IN_CHANX_N23751_37,IN_CHANX_N23750_36,IN_CHANX_N23749_29,
    IN_CHANX_N23748_28,IN_CHANX_N23747_21}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN23_N14785_io_in_hi = {IN_CHANX_N23771_7,IN_CHANX_N23770_6,IN_CHANX_N23755_53,IN_CHANX_N23754_52,
    IN_CHANX_N23753_45,IN_CHANX_N23752_44,CBMux_IPIN23_N14785_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN24_N14786_io_in_lo_lo = {IN_CHANX_N23756_60,_CBMux_IPIN19_N14781_io_in_WIRE_1,IN_CHANX_N23702_80,
    _CBMux_IPIN16_N14778_io_in_WIRE_1,IN_CHANX_N23682_0}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN24_N14786_io_in_lo = {IN_CHANX_N23772_14,IN_CHANX_N23761_77,IN_CHANX_N23760_76,
    IN_CHANX_N23759_69,IN_CHANX_N23758_68,IN_CHANX_N23757_61,CBMux_IPIN24_N14786_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN24_N14786_io_in_hi_lo = {IN_CHANX_N23777_31,IN_CHANX_N23776_30,IN_CHANX_N23775_23,
    IN_CHANX_N23774_22,IN_CHANX_N23773_15}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN24_N14786_io_in_hi = {IN_CHANX_N23783_55,IN_CHANX_N23782_54,IN_CHANX_N23781_47,
    IN_CHANX_N23780_46,IN_CHANX_N23779_39,IN_CHANX_N23778_38,CBMux_IPIN24_N14786_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN25_N14787_io_in_lo_lo = {IN_CHANX_N23688_24,_CBMux_IPIN16_N14778_io_in_WIRE_5,IN_CHANX_N23686_16,
    _CBMux_IPIN16_N14778_io_in_WIRE_3,IN_CHANX_N23684_8}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN25_N14787_io_in_lo = {IN_CHANX_N23694_48,_CBMux_IPIN17_N14779_io_in_WIRE_1,IN_CHANX_N23692_40,
    _CBMux_IPIN16_N14778_io_in_WIRE_9,IN_CHANX_N23690_32,_CBMux_IPIN16_N14778_io_in_WIRE_7,
    CBMux_IPIN25_N14787_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN25_N14787_io_in_hi_lo = {IN_CHANX_N23715_11,IN_CHANX_N23714_10,IN_CHANX_N23713_3,
    IN_CHANX_N23712_2,_CBMux_IPIN17_N14779_io_in_WIRE_3}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN25_N14787_io_in_hi = {IN_CHANX_N23789_79,IN_CHANX_N23788_78,IN_CHANX_N23787_71,
    IN_CHANX_N23786_70,IN_CHANX_N23785_63,IN_CHANX_N23784_62,CBMux_IPIN25_N14787_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN26_N14788_io_in_lo_lo = {_CBMux_IPIN17_N14779_io_in_WIRE_9,IN_CHANX_N23700_72,
    _CBMux_IPIN17_N14779_io_in_WIRE_7,IN_CHANX_N23698_64,_CBMux_IPIN17_N14779_io_in_WIRE_5,IN_CHANX_N23696_56}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN26_N14788_io_in_lo = {IN_CHANX_N23722_42,IN_CHANX_N23721_35,IN_CHANX_N23720_34,
    IN_CHANX_N23719_27,IN_CHANX_N23718_26,IN_CHANX_N23717_19,IN_CHANX_N23716_18,CBMux_IPIN26_N14788_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN26_N14788_io_in_hi_lo = {IN_CHANX_N23742_4,IN_CHANX_N23727_59,IN_CHANX_N23726_58,
    IN_CHANX_N23725_51,IN_CHANX_N23724_50,IN_CHANX_N23723_43}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN26_N14788_io_in_hi = {IN_CHANX_N23793_95,IN_CHANX_N23792_94,IN_CHANX_N23791_87,
    IN_CHANX_N23790_86,IN_CHANX_N23745_13,IN_CHANX_N23744_12,IN_CHANX_N23743_5,CBMux_IPIN26_N14788_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN27_N14789_io_in_lo_lo = {IN_CHANX_N23723_43,IN_CHANX_N23722_42,_CBMux_IPIN17_N14779_io_in_WIRE_13
    ,IN_CHANX_N23706_96,_CBMux_IPIN17_N14779_io_in_WIRE_11,IN_CHANX_N23704_88}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN27_N14789_io_in_lo = {IN_CHANX_N23730_74,IN_CHANX_N23729_67,IN_CHANX_N23728_66,
    IN_CHANX_N23727_59,IN_CHANX_N23726_58,IN_CHANX_N23725_51,IN_CHANX_N23724_50,CBMux_IPIN27_N14789_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN27_N14789_io_in_hi_lo = {IN_CHANX_N23744_12,IN_CHANX_N23743_5,IN_CHANX_N23742_4,
    IN_CHANX_N23733_83,IN_CHANX_N23732_82,IN_CHANX_N23731_75}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN27_N14789_io_in_hi = {IN_CHANX_N23751_37,IN_CHANX_N23750_36,IN_CHANX_N23749_29,
    IN_CHANX_N23748_28,IN_CHANX_N23747_21,IN_CHANX_N23746_20,IN_CHANX_N23745_13,CBMux_IPIN27_N14789_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN28_N14790_io_in_lo_lo = {IN_CHANX_N23729_67,IN_CHANX_N23728_66,_CBMux_IPIN17_N14779_io_in_WIRE_13
    ,IN_CHANX_N23706_96,_CBMux_IPIN17_N14779_io_in_WIRE_11,IN_CHANX_N23704_88}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN28_N14790_io_in_lo = {IN_CHANX_N23748_28,IN_CHANX_N23747_21,IN_CHANX_N23746_20,
    IN_CHANX_N23733_83,IN_CHANX_N23732_82,IN_CHANX_N23731_75,IN_CHANX_N23730_74,CBMux_IPIN28_N14790_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN28_N14790_io_in_hi_lo = {IN_CHANX_N23754_52,IN_CHANX_N23753_45,IN_CHANX_N23752_44,
    IN_CHANX_N23751_37,IN_CHANX_N23750_36,IN_CHANX_N23749_29}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN28_N14790_io_in_hi = {IN_CHANX_N23773_15,IN_CHANX_N23772_14,IN_CHANX_N23771_7,IN_CHANX_N23770_6,
    IN_CHANX_N23757_61,IN_CHANX_N23756_60,IN_CHANX_N23755_53,CBMux_IPIN28_N14790_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN29_N14791_io_in_lo_lo = {IN_CHANX_N23702_80,_CBMux_IPIN16_N14778_io_in_WIRE_3,IN_CHANX_N23684_8,
    _CBMux_IPIN16_N14778_io_in_WIRE_1,IN_CHANX_N23682_0}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN29_N14791_io_in_lo = {IN_CHANX_N23774_22,IN_CHANX_N23761_77,IN_CHANX_N23760_76,
    IN_CHANX_N23759_69,IN_CHANX_N23758_68,_CBMux_IPIN19_N14781_io_in_WIRE_1,CBMux_IPIN29_N14791_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN29_N14791_io_in_hi_lo = {IN_CHANX_N23779_39,IN_CHANX_N23778_38,IN_CHANX_N23777_31,
    IN_CHANX_N23776_30,IN_CHANX_N23775_23}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN29_N14791_io_in_hi = {IN_CHANX_N23785_63,IN_CHANX_N23784_62,IN_CHANX_N23783_55,
    IN_CHANX_N23782_54,IN_CHANX_N23781_47,IN_CHANX_N23780_46,CBMux_IPIN29_N14791_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN30_N14792_io_in_lo_lo = {IN_CHANX_N23690_32,_CBMux_IPIN16_N14778_io_in_WIRE_7,IN_CHANX_N23688_24,
    _CBMux_IPIN16_N14778_io_in_WIRE_5,IN_CHANX_N23686_16}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN30_N14792_io_in_lo = {IN_CHANX_N23696_56,_CBMux_IPIN17_N14779_io_in_WIRE_3,IN_CHANX_N23694_48,
    _CBMux_IPIN17_N14779_io_in_WIRE_1,IN_CHANX_N23692_40,_CBMux_IPIN16_N14778_io_in_WIRE_9,
    CBMux_IPIN30_N14792_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN30_N14792_io_in_hi_lo = {IN_CHANX_N23715_11,IN_CHANX_N23714_10,IN_CHANX_N23713_3,
    IN_CHANX_N23712_2,_CBMux_IPIN17_N14779_io_in_WIRE_5}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN30_N14792_io_in_hi = {IN_CHANX_N23789_79,IN_CHANX_N23788_78,IN_CHANX_N23787_71,
    IN_CHANX_N23786_70,IN_CHANX_N23717_19,IN_CHANX_N23716_18,CBMux_IPIN30_N14792_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN32_N14794_io_in_lo_lo = {IN_CHANX_N23733_83,IN_CHANX_N23732_82,IN_CHANX_N23731_75,
    IN_CHANX_N23730_74,IN_CHANX_N23729_67,IN_CHANX_N23728_66}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN32_N14794_io_in_lo = {IN_CHANX_N23752_44,IN_CHANX_N23751_37,IN_CHANX_N23750_36,
    IN_CHANX_N23749_29,IN_CHANX_N23748_28,IN_CHANX_N23747_21,IN_CHANX_N23746_20,CBMux_IPIN32_N14794_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN32_N14794_io_in_hi_lo = {IN_CHANX_N23770_6,IN_CHANX_N23757_61,IN_CHANX_N23756_60,
    IN_CHANX_N23755_53,IN_CHANX_N23754_52,IN_CHANX_N23753_45}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN32_N14794_io_in_hi = {IN_CHANX_N23793_95,IN_CHANX_N23792_94,IN_CHANX_N23791_87,
    IN_CHANX_N23790_86,IN_CHANX_N23773_15,IN_CHANX_N23772_14,IN_CHANX_N23771_7,CBMux_IPIN32_N14794_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN33_N14795_io_in_lo_lo = {_CBMux_IPIN19_N14781_io_in_WIRE_1,IN_CHANX_N23702_80,
    _CBMux_IPIN16_N14778_io_in_WIRE_3,IN_CHANX_N23684_8,_CBMux_IPIN16_N14778_io_in_WIRE_1,IN_CHANX_N23682_0}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN33_N14795_io_in_lo = {IN_CHANX_N23760_76,IN_CHANX_N23759_69,IN_CHANX_N23758_68,
    _CBMux_IPIN17_N14779_io_in_WIRE_13,IN_CHANX_N23706_96,_CBMux_IPIN17_N14779_io_in_WIRE_11,IN_CHANX_N23704_88,
    CBMux_IPIN33_N14795_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN33_N14795_io_in_hi_lo = {IN_CHANX_N23778_38,IN_CHANX_N23777_31,IN_CHANX_N23776_30,
    IN_CHANX_N23775_23,IN_CHANX_N23774_22,IN_CHANX_N23761_77}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN33_N14795_io_in_hi = {IN_CHANX_N23785_63,IN_CHANX_N23784_62,IN_CHANX_N23783_55,
    IN_CHANX_N23782_54,IN_CHANX_N23781_47,IN_CHANX_N23780_46,IN_CHANX_N23779_39,CBMux_IPIN33_N14795_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN35_N14797_io_in_lo_lo = {IN_CHANX_N23694_48,_CBMux_IPIN17_N14779_io_in_WIRE_1,IN_CHANX_N23692_40,
    _CBMux_IPIN16_N14778_io_in_WIRE_9,IN_CHANX_N23690_32}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN35_N14797_io_in_lo = {IN_CHANX_N23700_72,_CBMux_IPIN17_N14779_io_in_WIRE_7,IN_CHANX_N23698_64,
    _CBMux_IPIN17_N14779_io_in_WIRE_5,IN_CHANX_N23696_56,_CBMux_IPIN17_N14779_io_in_WIRE_3,
    CBMux_IPIN35_N14797_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN35_N14797_io_in_hi_lo = {IN_CHANX_N23715_11,IN_CHANX_N23714_10,IN_CHANX_N23713_3,
    IN_CHANX_N23712_2,_CBMux_IPIN17_N14779_io_in_WIRE_9}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN35_N14797_io_in_hi = {IN_CHANX_N23721_35,IN_CHANX_N23720_34,IN_CHANX_N23719_27,
    IN_CHANX_N23718_26,IN_CHANX_N23717_19,IN_CHANX_N23716_18,CBMux_IPIN35_N14797_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN36_N14798_io_in_lo = {IN_CHANX_N23748_28,IN_CHANX_N23747_21,IN_CHANX_N23746_20,
    IN_CHANX_N23733_83,IN_CHANX_N23732_82,IN_CHANX_N23731_75,CBMux_IPIN23_N14785_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN36_N14798_io_in_hi_lo = {IN_CHANX_N23753_45,IN_CHANX_N23752_44,IN_CHANX_N23751_37,
    IN_CHANX_N23750_36,IN_CHANX_N23749_29}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN36_N14798_io_in_hi = {IN_CHANX_N23773_15,IN_CHANX_N23772_14,IN_CHANX_N23771_7,IN_CHANX_N23770_6,
    IN_CHANX_N23755_53,IN_CHANX_N23754_52,CBMux_IPIN36_N14798_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN37_N14799_io_in_lo_lo = {IN_CHANX_N23757_61,IN_CHANX_N23756_60,_CBMux_IPIN19_N14781_io_in_WIRE_1,
    IN_CHANX_N23702_80,_CBMux_IPIN16_N14778_io_in_WIRE_1,IN_CHANX_N23682_0}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN37_N14799_io_in_lo = {IN_CHANX_N23774_22,IN_CHANX_N23773_15,IN_CHANX_N23772_14,
    IN_CHANX_N23761_77,IN_CHANX_N23760_76,IN_CHANX_N23759_69,IN_CHANX_N23758_68,CBMux_IPIN37_N14799_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN37_N14799_io_in_hi_lo = {IN_CHANX_N23780_46,IN_CHANX_N23779_39,IN_CHANX_N23778_38,
    IN_CHANX_N23777_31,IN_CHANX_N23776_30,IN_CHANX_N23775_23}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN37_N14799_io_in_hi = {IN_CHANX_N23793_95,IN_CHANX_N23792_94,IN_CHANX_N23791_87,
    IN_CHANX_N23790_86,IN_CHANX_N23783_55,IN_CHANX_N23782_54,IN_CHANX_N23781_47,CBMux_IPIN37_N14799_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN38_N14800_io_in_lo = {IN_CHANX_N23714_10,_CBMux_IPIN17_N14779_io_in_WIRE_13,IN_CHANX_N23706_96,
    _CBMux_IPIN17_N14779_io_in_WIRE_11,IN_CHANX_N23704_88,_CBMux_IPIN17_N14779_io_in_WIRE_9,IN_CHANX_N23700_72,
    CBMux_IPIN22_N14784_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [5:0] CBMux_IPIN38_N14800_io_in_hi_lo = {IN_CHANX_N23720_34,IN_CHANX_N23719_27,IN_CHANX_N23718_26,
    IN_CHANX_N23717_19,IN_CHANX_N23716_18,IN_CHANX_N23715_11}; // @[TileFull.scala 175:8]
  wire [12:0] CBMux_IPIN38_N14800_io_in_hi = {IN_CHANX_N23743_5,IN_CHANX_N23742_4,IN_CHANX_N23725_51,IN_CHANX_N23724_50,
    IN_CHANX_N23723_43,IN_CHANX_N23722_42,IN_CHANX_N23721_35,CBMux_IPIN38_N14800_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN39_N14801_io_in_lo_lo = {IN_CHANX_N23686_16,_CBMux_IPIN16_N14778_io_in_WIRE_3,IN_CHANX_N23684_8,
    _CBMux_IPIN16_N14778_io_in_WIRE_1,IN_CHANX_N23682_0}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN39_N14801_io_in_lo = {IN_CHANX_N23778_38,_CBMux_IPIN19_N14781_io_in_WIRE_1,IN_CHANX_N23702_80,
    _CBMux_IPIN16_N14778_io_in_WIRE_7,IN_CHANX_N23688_24,_CBMux_IPIN16_N14778_io_in_WIRE_5,
    CBMux_IPIN39_N14801_io_in_lo_lo}; // @[TileFull.scala 175:8]
  wire [4:0] CBMux_IPIN39_N14801_io_in_hi_lo = {IN_CHANX_N23783_55,IN_CHANX_N23782_54,IN_CHANX_N23781_47,
    IN_CHANX_N23780_46,IN_CHANX_N23779_39}; // @[TileFull.scala 175:8]
  wire [10:0] CBMux_IPIN39_N14801_io_in_hi = {IN_CHANX_N23789_79,IN_CHANX_N23788_78,IN_CHANX_N23787_71,
    IN_CHANX_N23786_70,IN_CHANX_N23785_63,IN_CHANX_N23784_62,CBMux_IPIN39_N14801_io_in_hi_lo}; // @[TileFull.scala 175:8]
  wire  _SBMux_C1_N23683_O_3_C_6_io_in_WIRE_1 = logicBlock_OPIN_83; // @[TileFull.scala 187:{39,39}]
  wire  _SBMux_C1_N23683_O_3_C_6_io_in_WIRE_0 = logicBlock_OPIN_81; // @[TileFull.scala 187:{39,39}]
  wire  _SBMux_C1_N23683_O_3_C_6_io_in_WIRE_2 = logicBlock_OPIN_86; // @[TileFull.scala 187:{39,39}]
  wire [3:0] SBMux_C1_N23683_O_3_C_6_io_in_lo = {IN_CHANY_N30094_16,_SBMux_C1_N23683_O_3_C_6_io_in_WIRE_2,
    _SBMux_C1_N23683_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N23683_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C1_N23683_O_3_C_6_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30211_97,IN_CHANY_N30178_100,
    IN_CHANY_N30166_88,IN_CHANY_N30149_71}; // @[TileFull.scala 202:13]
  wire  _SBMux_C9_N23685_O_3_C_7_io_in_WIRE_1 = logicBlock_OPIN_84; // @[TileFull.scala 187:{39,39}]
  wire [4:0] SBMux_C9_N23685_O_3_C_7_io_in_lo = {IN_CHANY_N30174_96,IN_CHANY_N30152_74,
    _SBMux_C1_N23683_O_3_C_6_io_in_WIRE_2,_SBMux_C9_N23685_O_3_C_7_io_in_WIRE_1,_SBMux_C1_N23683_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C9_N23685_O_3_C_7_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30213_101,IN_CHANY_N30211_97,
    IN_CHANY_N30195_33,IN_CHANY_N30182_104}; // @[TileFull.scala 202:13]
  wire  _SBMux_C17_N23687_O_3_C_6_io_in_WIRE_2 = logicBlock_OPIN_87; // @[TileFull.scala 187:{39,39}]
  wire [3:0] SBMux_C17_N23687_O_3_C_6_io_in_lo = {IN_CHANY_N30092_14,_SBMux_C17_N23687_O_3_C_6_io_in_WIRE_2,
    _SBMux_C9_N23685_O_3_C_7_io_in_WIRE_1,_SBMux_C1_N23683_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C17_N23687_O_3_C_6_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30211_97,IN_CHANY_N30178_100,
    IN_CHANY_N30166_88,IN_CHANY_N30141_63}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C25_N23689_O_3_C_6_io_in_lo = {IN_CHANY_N30107_29,_SBMux_C17_N23687_O_3_C_6_io_in_WIRE_2,
    _SBMux_C9_N23685_O_3_C_7_io_in_WIRE_1,_SBMux_C1_N23683_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C25_N23689_O_3_C_6_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30209_89,IN_CHANY_N30182_104,
    IN_CHANY_N30174_96,IN_CHANY_N30138_60}; // @[TileFull.scala 202:13]
  wire  _SBMux_C33_N23691_O_3_C_7_io_in_WIRE_0 = logicBlock_OPIN_82; // @[TileFull.scala 187:{39,39}]
  wire [4:0] SBMux_C33_N23691_O_3_C_7_io_in_lo = {IN_CHANY_N30160_82,IN_CHANY_N30113_35,
    _SBMux_C17_N23687_O_3_C_6_io_in_WIRE_2,_SBMux_C9_N23685_O_3_C_7_io_in_WIRE_1,_SBMux_C33_N23691_O_3_C_7_io_in_WIRE_0}
    ; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C33_N23691_O_3_C_7_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30211_97,IN_CHANY_N30209_89,
    IN_CHANY_N30178_100,IN_CHANY_N30174_96}; // @[TileFull.scala 202:13]
  wire  _SBMux_C41_N23693_O_3_C_6_io_in_WIRE_1 = logicBlock_OPIN_85; // @[TileFull.scala 187:{39,39}]
  wire [3:0] SBMux_C41_N23693_O_3_C_6_io_in_lo = {IN_CHANY_N30080_2,_SBMux_C17_N23687_O_3_C_6_io_in_WIRE_2,
    _SBMux_C41_N23693_O_3_C_6_io_in_WIRE_1,_SBMux_C33_N23691_O_3_C_7_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C41_N23693_O_3_C_6_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30209_89,IN_CHANY_N30178_100,
    IN_CHANY_N30174_96,IN_CHANY_N30133_55}; // @[TileFull.scala 202:13]
  wire  _SBMux_C49_N23695_O_3_C_5_io_in_WIRE_2 = logicBlock_OPIN_88; // @[TileFull.scala 187:{39,39}]
  wire [3:0] SBMux_C49_N23695_O_3_C_5_io_in_lo = {IN_CHANY_N30109_31,_SBMux_C49_N23695_O_3_C_5_io_in_WIRE_2,
    _SBMux_C41_N23693_O_3_C_6_io_in_WIRE_1,_SBMux_C33_N23691_O_3_C_7_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C49_N23695_O_3_C_5_io_in_hi = {IN_CHANY_N30211_97,IN_CHANY_N30182_104,IN_CHANY_N30166_88,
    IN_CHANY_N30114_36}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C57_N23697_O_3_C_6_io_in_lo = {IN_CHANY_N30105_27,_SBMux_C49_N23695_O_3_C_5_io_in_WIRE_2,
    _SBMux_C41_N23693_O_3_C_6_io_in_WIRE_1,_SBMux_C33_N23691_O_3_C_7_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C57_N23697_O_3_C_6_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30209_89,IN_CHANY_N30178_100,
    IN_CHANY_N30166_88,IN_CHANY_N30120_42}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C65_N23699_O_3_C_6_io_in_lo = {IN_CHANY_N30098_20,_SBMux_C49_N23695_O_3_C_5_io_in_WIRE_2,
    _SBMux_C41_N23693_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N23683_O_3_C_6_io_in_WIRE_1}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C65_N23699_O_3_C_6_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30209_89,IN_CHANY_N30193_25,
    IN_CHANY_N30182_104,IN_CHANY_N30166_88}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C73_N23701_O_3_C_6_io_in_lo = {IN_CHANY_N30100_22,_SBMux_C49_N23695_O_3_C_5_io_in_WIRE_2,
    _SBMux_C1_N23683_O_3_C_6_io_in_WIRE_2,_SBMux_C1_N23683_O_3_C_6_io_in_WIRE_1}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C73_N23701_O_3_C_6_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30211_97,IN_CHANY_N30178_100,
    IN_CHANY_N30166_88,IN_CHANY_N30145_67}; // @[TileFull.scala 202:13]
  wire [2:0] SBMux_C81_N23703_O_2_C_5_io_in_lo = {IN_CHANY_N30088_10,_SBMux_C1_N23683_O_3_C_6_io_in_WIRE_2,
    _SBMux_C1_N23683_O_3_C_6_io_in_WIRE_1}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C81_N23703_O_2_C_5_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30182_104,IN_CHANY_N30174_96,
    IN_CHANY_N30153_75}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C89_N23705_O_3_C_5_io_in_lo = {IN_CHANX_N23821_89,_SBMux_C41_N23693_O_3_C_6_io_in_WIRE_1,
    _SBMux_C1_N23683_O_3_C_6_io_in_WIRE_1,_SBMux_C1_N23683_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C89_N23705_O_3_C_5_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30209_89,IN_CHANY_N30182_104,
    IN_CHANY_N30174_96}; // @[TileFull.scala 202:13]
  wire [2:0] SBMux_C97_N23707_O_2_C_5_io_in_lo = {IN_CHANX_N23823_97,_SBMux_C9_N23685_O_3_C_7_io_in_WIRE_1,
    _SBMux_C33_N23691_O_3_C_7_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C97_N23707_O_2_C_5_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30211_97,IN_CHANY_N30178_100,
    IN_CHANY_N30166_88}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C0_N23798_O_3_C_6_io_in_lo = {IN_CHANY_N30083_5,IN_OPIN_N17288_86,IN_OPIN_N17285_83,IN_OPIN_N17283_81
    }; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C0_N23798_O_3_C_6_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30209_89,IN_CHANY_N30178_100,
    IN_CHANY_N30166_88,IN_CHANY_N30156_78}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C8_N23800_O_3_C_6_io_in_lo = {IN_CHANY_N30150_72,IN_OPIN_N17288_86,IN_OPIN_N17286_84,
    IN_OPIN_N17283_81}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C8_N23800_O_3_C_6_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30209_89,IN_CHANY_N30205_73,
    IN_CHANY_N30182_104,IN_CHANY_N30174_96}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C16_N23802_O_3_C_6_io_in_lo = {IN_CHANY_N30104_26,IN_OPIN_N17289_87,IN_OPIN_N17286_84,
    IN_OPIN_N17283_81}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C16_N23802_O_3_C_6_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30209_89,IN_CHANY_N30182_104,
    IN_CHANY_N30174_96,IN_CHANY_N30137_59}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C24_N23804_O_3_C_7_io_in_lo = {IN_CHANY_N30149_71,IN_CHANY_N30130_52,IN_OPIN_N17289_87,
    IN_OPIN_N17286_84,IN_OPIN_N17283_81}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C24_N23804_O_3_C_7_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30209_89,IN_CHANY_N30182_104,
    IN_CHANY_N30178_100,IN_CHANY_N30166_88}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C32_N23806_O_3_C_5_io_in_lo = {IN_CHANY_N30136_58,IN_OPIN_N17289_87,IN_OPIN_N17286_84,
    IN_OPIN_N17284_82}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C32_N23806_O_3_C_5_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30211_97,IN_CHANY_N30201_57,
    IN_CHANY_N30182_104}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C40_N23808_O_3_C_5_io_in_lo = {IN_CHANY_N30118_40,IN_OPIN_N17289_87,IN_OPIN_N17287_85,
    IN_OPIN_N17284_82}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C40_N23808_O_3_C_5_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30211_97,IN_CHANY_N30199_49,
    IN_CHANY_N30174_96}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C48_N23810_O_3_C_6_io_in_lo = {IN_CHANY_N30081_3,IN_OPIN_N17290_88,IN_OPIN_N17287_85,
    IN_OPIN_N17284_82}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C48_N23810_O_3_C_6_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30211_97,IN_CHANY_N30178_100,
    IN_CHANY_N30174_96,IN_CHANY_N30116_38}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C56_N23812_O_3_C_6_io_in_lo = {IN_CHANY_N30123_45,IN_OPIN_N17290_88,IN_OPIN_N17287_85,
    IN_OPIN_N17284_82}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C56_N23812_O_3_C_6_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30209_89,IN_CHANY_N30182_104,
    IN_CHANY_N30166_88,IN_CHANY_N30158_80}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C64_N23814_O_3_C_6_io_in_lo = {IN_CHANY_N30084_6,IN_OPIN_N17290_88,IN_OPIN_N17287_85,
    IN_OPIN_N17285_83}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C64_N23814_O_3_C_6_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30211_97,IN_CHANY_N30178_100,
    IN_CHANY_N30166_88,IN_CHANY_N30109_31}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C72_N23816_O_3_C_7_io_in_lo = {IN_CHANY_N30134_56,IN_CHANY_N30101_23,IN_OPIN_N17290_88,
    IN_OPIN_N17288_86,IN_OPIN_N17285_83}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C72_N23816_O_3_C_7_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30211_97,IN_CHANY_N30178_100,
    IN_CHANY_N30174_96,IN_CHANY_N30166_88}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C80_N23818_O_2_C_6_io_in_lo = {IN_CHANY_N30141_63,IN_CHANY_N30102_24,IN_OPIN_N17288_86,
    IN_OPIN_N17285_83}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C80_N23818_O_2_C_6_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30211_97,IN_CHANY_N30182_104,
    IN_CHANY_N30166_88}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C88_N23820_O_3_C_5_io_in_lo = {IN_CHANX_N23704_88,IN_OPIN_N17287_85,IN_OPIN_N17285_83,
    IN_OPIN_N17283_81}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C88_N23820_O_3_C_5_io_in_hi = {IN_CHANY_N30215_105,IN_CHANY_N30211_97,IN_CHANY_N30182_104,
    IN_CHANY_N30174_96}; // @[TileFull.scala 202:13]
  wire [2:0] SBMux_C96_N23822_O_2_C_5_io_in_lo = {IN_CHANX_N23706_96,IN_OPIN_N17286_84,IN_OPIN_N17284_82}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C96_N23822_O_2_C_5_io_in_hi = {IN_CHANY_N30213_101,IN_CHANY_N30209_89,IN_CHANY_N30178_100,
    IN_CHANY_N30166_88}; // @[TileFull.scala 202:13]
  wire  _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_1 = logicBlock_OPIN_75; // @[TileFull.scala 187:{39,39}]
  wire  _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_0 = logicBlock_OPIN_73; // @[TileFull.scala 187:{39,39}]
  wire [1:0] SBMux_C1_N30079_O_4_C_6_io_in_lo_lo = {_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_1,
    _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire  _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_3 = logicBlock_OPIN_80; // @[TileFull.scala 187:{39,39}]
  wire  _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_2 = logicBlock_OPIN_77; // @[TileFull.scala 187:{39,39}]
  wire [4:0] SBMux_C1_N30079_O_4_C_6_io_in_lo = {IN_CHANX_N23704_88,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_3,
    _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_2,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_1,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C1_N30079_O_4_C_6_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23823_97,IN_CHANX_N23766_100,
    IN_CHANX_N23748_28,IN_CHANX_N23745_13}; // @[TileFull.scala 202:13]
  wire  _SBMux_C9_N30087_O_4_C_7_io_in_WIRE_2 = logicBlock_OPIN_78; // @[TileFull.scala 187:{39,39}]
  wire [4:0] SBMux_C9_N30087_O_4_C_7_io_in_lo = {IN_CHANX_N23704_88,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_3,
    _SBMux_C9_N30087_O_4_C_7_io_in_WIRE_2,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_1,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [5:0] SBMux_C9_N30087_O_4_C_7_io_in_hi = {IN_CHANX_N23827_105,IN_CHANX_N23823_97,IN_CHANX_N23821_89,
    IN_CHANX_N23777_31,IN_CHANX_N23766_100,IN_CHANX_N23742_4}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C17_N30095_O_3_C_7_io_in_lo = {IN_CHANX_N23704_88,IN_CHANX_N23700_72,
    _SBMux_C9_N30087_O_4_C_7_io_in_WIRE_2,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_1,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C17_N30095_O_3_C_7_io_in_hi = {IN_CHANX_N23827_105,IN_CHANX_N23825_101,IN_CHANX_N23821_89,
    IN_CHANX_N23799_1,IN_CHANX_N23768_104}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C25_N30103_O_3_C_6_io_in_lo = {IN_CHANX_N23704_88,_SBMux_C9_N30087_O_4_C_7_io_in_WIRE_2,
    _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_1,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C25_N30103_O_3_C_6_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23821_89,IN_CHANX_N23766_100,
    IN_CHANX_N23728_66,IN_CHANX_N23713_3}; // @[TileFull.scala 202:13]
  wire  _SBMux_C33_N30111_O_3_C_4_io_in_WIRE_1 = logicBlock_OPIN_76; // @[TileFull.scala 187:{39,39}]
  wire [2:0] SBMux_C33_N30111_O_3_C_4_io_in_lo = {_SBMux_C9_N30087_O_4_C_7_io_in_WIRE_2,
    _SBMux_C33_N30111_O_3_C_4_io_in_WIRE_1,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C33_N30111_O_3_C_4_io_in_hi = {IN_CHANX_N23766_100,IN_CHANX_N23723_43,IN_CHANX_N23704_88,
    IN_CHANX_N23690_32}; // @[TileFull.scala 202:13]
  wire  _SBMux_C41_N30119_O_3_C_6_io_in_WIRE_0 = logicBlock_OPIN_74; // @[TileFull.scala 187:{39,39}]
  wire [1:0] SBMux_C41_N30119_O_3_C_6_io_in_lo_lo = {_SBMux_C33_N30111_O_3_C_4_io_in_WIRE_1,
    _SBMux_C41_N30119_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire  _SBMux_C41_N30119_O_3_C_6_io_in_WIRE_2 = logicBlock_OPIN_79; // @[TileFull.scala 187:{39,39}]
  wire [3:0] SBMux_C41_N30119_O_3_C_6_io_in_lo = {IN_CHANX_N23706_96,_SBMux_C41_N30119_O_3_C_6_io_in_WIRE_2,
    _SBMux_C33_N30111_O_3_C_4_io_in_WIRE_1,_SBMux_C41_N30119_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C41_N30119_O_3_C_6_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23821_89,IN_CHANX_N23782_54,
    IN_CHANX_N23766_100,IN_CHANX_N23753_45}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C49_N30127_O_3_C_6_io_in_hi = {IN_CHANX_N23827_105,IN_CHANX_N23823_97,IN_CHANX_N23801_9,
    IN_CHANX_N23768_104,IN_CHANX_N23744_12}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C57_N30135_O_3_C_6_io_in_lo = {IN_CHANX_N23692_40,_SBMux_C41_N30119_O_3_C_6_io_in_WIRE_2,
    _SBMux_C33_N30111_O_3_C_4_io_in_WIRE_1,_SBMux_C41_N30119_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C57_N30135_O_3_C_6_io_in_hi = {IN_CHANX_N23827_105,IN_CHANX_N23823_97,IN_CHANX_N23781_47,
    IN_CHANX_N23768_104,IN_CHANX_N23704_88}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C65_N30143_O_3_C_6_io_in_lo = {IN_CHANX_N23706_96,_SBMux_C41_N30119_O_3_C_6_io_in_WIRE_2,
    _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_2,_SBMux_C41_N30119_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C65_N30143_O_3_C_6_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23821_89,IN_CHANX_N23813_57,
    IN_CHANX_N23768_104,IN_CHANX_N23730_74}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C73_N30151_O_3_C_6_io_in_lo = {IN_CHANX_N23706_96,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_3,
    _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_2,_SBMux_C41_N30119_O_3_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C73_N30151_O_3_C_6_io_in_hi = {IN_CHANX_N23827_105,IN_CHANX_N23821_89,IN_CHANX_N23778_38,
    IN_CHANX_N23766_100,IN_CHANX_N23759_69}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C81_N30159_O_3_C_6_io_in_lo = {IN_CHANX_N23706_96,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_3,
    _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_2,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_1}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C81_N30159_O_3_C_6_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23823_97,IN_CHANX_N23775_23,
    IN_CHANX_N23768_104,IN_CHANX_N23718_26}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C89_N30167_O_4_C_5_io_in_lo = {_SBMux_C41_N30119_O_3_C_6_io_in_WIRE_2,
    _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_2,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_1,_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_0}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C89_N30167_O_4_C_5_io_in_hi = {IN_CHANY_N30209_89,IN_CHANX_N23827_105,IN_CHANX_N23823_97,
    IN_CHANX_N23766_100,IN_CHANX_N23706_96}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C97_N30175_O_4_C_5_io_in_lo = {_SBMux_C1_N30079_O_4_C_6_io_in_WIRE_3,
    _SBMux_C9_N30087_O_4_C_7_io_in_WIRE_2,_SBMux_C33_N30111_O_3_C_4_io_in_WIRE_1,_SBMux_C41_N30119_O_3_C_6_io_in_WIRE_0}
    ; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C97_N30175_O_4_C_5_io_in_hi = {IN_CHANY_N30211_97,IN_CHANX_N23825_101,IN_CHANX_N23821_89,
    IN_CHANX_N23768_104,IN_CHANX_N23704_88}; // @[TileFull.scala 202:13]
  wire [2:0] SBMux_C101_N30179_O_4_C_1_io_in_hi = {IN_CHANY_N30215_105,_SBMux_C41_N30119_O_3_C_6_io_in_WIRE_2,
    _SBMux_C1_N30079_O_4_C_6_io_in_WIRE_2}; // @[TileFull.scala 202:13]
  wire [1:0] SBMux_C105_N30183_O_3_C_1_io_in_hi = {IN_CHANY_N30213_101,_SBMux_C9_N30087_O_4_C_7_io_in_WIRE_2}; // @[TileFull.scala 202:13]
  wire [1:0] SBMux_C0_N30186_O_4_C_6_io_in_lo_lo = {IN_OPIN_N15081_75,IN_OPIN_N15079_73}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C0_N30186_O_4_C_6_io_in_lo = {IN_CHANX_N23688_24,IN_OPIN_N15086_80,IN_OPIN_N15083_77,
    IN_OPIN_N15081_75,IN_OPIN_N15079_73}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C0_N30186_O_4_C_6_io_in_hi = {IN_CHANX_N23827_105,IN_CHANX_N23823_97,IN_CHANX_N23768_104,
    IN_CHANX_N23761_77,IN_CHANX_N23704_88}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C8_N30188_O_4_C_5_io_in_lo = {IN_OPIN_N15086_80,IN_OPIN_N15084_78,IN_OPIN_N15081_75,IN_OPIN_N15079_73
    }; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C8_N30188_O_4_C_5_io_in_hi = {IN_CHANX_N23827_105,IN_CHANX_N23821_89,IN_CHANX_N23809_41,
    IN_CHANX_N23766_100,IN_CHANX_N23742_4}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C16_N30190_O_3_C_7_io_in_lo = {IN_CHANX_N23706_96,IN_CHANX_N23704_88,IN_OPIN_N15084_78,
    IN_OPIN_N15081_75,IN_OPIN_N15079_73}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C16_N30190_O_3_C_7_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23823_97,IN_CHANX_N23781_47,
    IN_CHANX_N23776_30,IN_CHANX_N23768_104}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C24_N30192_O_3_C_6_io_in_lo = {IN_CHANX_N23704_88,IN_OPIN_N15084_78,IN_OPIN_N15081_75,
    IN_OPIN_N15079_73}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C24_N30192_O_3_C_6_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23823_97,IN_CHANX_N23803_17,
    IN_CHANX_N23766_100,IN_CHANX_N23718_26}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C32_N30194_O_3_C_6_io_in_lo = {IN_CHANX_N23704_88,IN_OPIN_N15084_78,IN_OPIN_N15082_76,
    IN_OPIN_N15079_73}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C32_N30194_O_3_C_6_io_in_hi = {IN_CHANX_N23827_105,IN_CHANX_N23823_97,IN_CHANX_N23770_6,
    IN_CHANX_N23768_104,IN_CHANX_N23729_67}; // @[TileFull.scala 202:13]
  wire [1:0] SBMux_C40_N30196_O_3_C_5_io_in_lo_lo = {IN_OPIN_N15082_76,IN_OPIN_N15080_74}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C40_N30196_O_3_C_5_io_in_lo = {IN_CHANX_N23706_96,IN_OPIN_N15085_79,IN_OPIN_N15082_76,
    IN_OPIN_N15080_74}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C40_N30196_O_3_C_5_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23823_97,IN_CHANX_N23747_21,
    IN_CHANX_N23744_12}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C48_N30198_O_3_C_6_io_in_lo = {IN_CHANX_N23684_8,IN_OPIN_N15085_79,IN_OPIN_N15082_76,
    IN_OPIN_N15080_74}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C48_N30198_O_3_C_6_io_in_hi = {IN_CHANX_N23827_105,IN_CHANX_N23821_89,IN_CHANX_N23766_100,
    IN_CHANX_N23745_13,IN_CHANX_N23706_96}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C56_N30200_O_3_C_6_io_in_lo = {IN_CHANX_N23700_72,IN_OPIN_N15085_79,IN_OPIN_N15082_76,
    IN_OPIN_N15080_74}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C56_N30200_O_3_C_6_io_in_hi = {IN_CHANX_N23827_105,IN_CHANX_N23821_89,IN_CHANX_N23766_100,
    IN_CHANX_N23731_75,IN_CHANX_N23706_96}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C64_N30202_O_3_C_7_io_in_lo = {IN_CHANX_N23712_2,IN_CHANX_N23704_88,IN_OPIN_N15085_79,
    IN_OPIN_N15083_77,IN_OPIN_N15080_74}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C64_N30202_O_3_C_7_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23823_97,IN_CHANX_N23768_104,
    IN_CHANX_N23766_100,IN_CHANX_N23719_27}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C72_N30204_O_3_C_6_io_in_lo = {IN_CHANX_N23706_96,IN_OPIN_N15086_80,IN_OPIN_N15083_77,
    IN_OPIN_N15080_74}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C72_N30204_O_3_C_6_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23821_89,IN_CHANX_N23780_46,
    IN_CHANX_N23768_104,IN_CHANX_N23757_61}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C80_N30206_O_3_C_6_io_in_lo = {IN_CHANX_N23706_96,IN_OPIN_N15086_80,IN_OPIN_N15083_77,
    IN_OPIN_N15081_75}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C80_N30206_O_3_C_6_io_in_hi = {IN_CHANX_N23825_101,IN_CHANX_N23821_89,IN_CHANX_N23773_15,
    IN_CHANX_N23768_104,IN_CHANX_N23730_74}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C88_N30208_O_4_C_5_io_in_lo = {IN_OPIN_N15085_79,IN_OPIN_N15083_77,IN_OPIN_N15081_75,
    IN_OPIN_N15079_73}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C88_N30208_O_4_C_5_io_in_hi = {IN_CHANY_N30166_88,IN_CHANX_N23827_105,IN_CHANX_N23823_97,
    IN_CHANX_N23766_100,IN_CHANX_N23706_96}; // @[TileFull.scala 202:13]
  wire [3:0] SBMux_C96_N30210_O_4_C_5_io_in_lo = {IN_OPIN_N15086_80,IN_OPIN_N15084_78,IN_OPIN_N15082_76,
    IN_OPIN_N15080_74}; // @[TileFull.scala 202:13]
  wire [4:0] SBMux_C96_N30210_O_4_C_5_io_in_hi = {IN_CHANY_N30174_96,IN_CHANX_N23825_101,IN_CHANX_N23821_89,
    IN_CHANX_N23768_104,IN_CHANX_N23704_88}; // @[TileFull.scala 202:13]
  wire [2:0] SBMux_C100_N30212_O_4_C_1_io_in_hi = {IN_CHANY_N30178_100,IN_OPIN_N15085_79,IN_OPIN_N15083_77}; // @[TileFull.scala 202:13]
  wire [1:0] SBMux_C104_N30214_O_3_C_1_io_in_hi = {IN_CHANY_N30182_104,IN_OPIN_N15084_78}; // @[TileFull.scala 202:13]
  CLBlut4N10Mul logicBlock ( // @[TileFull.scala 47:37]
    .IPIN_0(logicBlock_IPIN_0),
    .IPIN_1(logicBlock_IPIN_1),
    .IPIN_2(logicBlock_IPIN_2),
    .IPIN_3(logicBlock_IPIN_3),
    .IPIN_4(logicBlock_IPIN_4),
    .IPIN_5(logicBlock_IPIN_5),
    .IPIN_6(logicBlock_IPIN_6),
    .IPIN_7(logicBlock_IPIN_7),
    .IPIN_8(logicBlock_IPIN_8),
    .IPIN_9(logicBlock_IPIN_9),
    .IPIN_10(logicBlock_IPIN_10),
    .IPIN_11(logicBlock_IPIN_11),
    .IPIN_12(logicBlock_IPIN_12),
    .IPIN_13(logicBlock_IPIN_13),
    .IPIN_14(logicBlock_IPIN_14),
    .IPIN_15(logicBlock_IPIN_15),
    .IPIN_16(logicBlock_IPIN_16),
    .IPIN_17(logicBlock_IPIN_17),
    .IPIN_18(logicBlock_IPIN_18),
    .IPIN_19(logicBlock_IPIN_19),
    .IPIN_20(logicBlock_IPIN_20),
    .IPIN_21(logicBlock_IPIN_21),
    .IPIN_22(logicBlock_IPIN_22),
    .IPIN_23(logicBlock_IPIN_23),
    .IPIN_24(logicBlock_IPIN_24),
    .IPIN_25(logicBlock_IPIN_25),
    .IPIN_26(logicBlock_IPIN_26),
    .IPIN_27(logicBlock_IPIN_27),
    .IPIN_28(logicBlock_IPIN_28),
    .IPIN_29(logicBlock_IPIN_29),
    .IPIN_30(logicBlock_IPIN_30),
    .IPIN_31(logicBlock_IPIN_31),
    .IPIN_32(logicBlock_IPIN_32),
    .IPIN_33(logicBlock_IPIN_33),
    .IPIN_34(logicBlock_IPIN_34),
    .IPIN_35(logicBlock_IPIN_35),
    .IPIN_36(logicBlock_IPIN_36),
    .IPIN_37(logicBlock_IPIN_37),
    .IPIN_38(logicBlock_IPIN_38),
    .IPIN_39(logicBlock_IPIN_39),
    .IPIN_40(logicBlock_IPIN_40),
    .IPIN_41(logicBlock_IPIN_41),
    .IPIN_42(logicBlock_IPIN_42),
    .IPIN_43(logicBlock_IPIN_43),
    .IPIN_44(logicBlock_IPIN_44),
    .IPIN_45(logicBlock_IPIN_45),
    .IPIN_46(logicBlock_IPIN_46),
    .IPIN_47(logicBlock_IPIN_47),
    .IPIN_48(logicBlock_IPIN_48),
    .IPIN_49(logicBlock_IPIN_49),
    .IPIN_50(logicBlock_IPIN_50),
    .IPIN_51(logicBlock_IPIN_51),
    .IPIN_52(logicBlock_IPIN_52),
    .IPIN_53(logicBlock_IPIN_53),
    .IPIN_54(logicBlock_IPIN_54),
    .IPIN_55(logicBlock_IPIN_55),
    .IPIN_56(logicBlock_IPIN_56),
    .IPIN_57(logicBlock_IPIN_57),
    .IPIN_58(logicBlock_IPIN_58),
    .IPIN_59(logicBlock_IPIN_59),
    .IPIN_60(logicBlock_IPIN_60),
    .IPIN_61(logicBlock_IPIN_61),
    .IPIN_62(logicBlock_IPIN_62),
    .IPIN_63(logicBlock_IPIN_63),
    .IPIN_64(logicBlock_IPIN_64),
    .IPIN_65(logicBlock_IPIN_65),
    .IPIN_66(logicBlock_IPIN_66),
    .IPIN_67(logicBlock_IPIN_67),
    .IPIN_68(logicBlock_IPIN_68),
    .IPIN_69(logicBlock_IPIN_69),
    .IPIN_70(logicBlock_IPIN_70),
    .IPIN_71(logicBlock_IPIN_71),
    .OPIN_73(logicBlock_OPIN_73),
    .OPIN_74(logicBlock_OPIN_74),
    .OPIN_75(logicBlock_OPIN_75),
    .OPIN_76(logicBlock_OPIN_76),
    .OPIN_77(logicBlock_OPIN_77),
    .OPIN_78(logicBlock_OPIN_78),
    .OPIN_79(logicBlock_OPIN_79),
    .OPIN_80(logicBlock_OPIN_80),
    .OPIN_81(logicBlock_OPIN_81),
    .OPIN_82(logicBlock_OPIN_82),
    .OPIN_83(logicBlock_OPIN_83),
    .OPIN_84(logicBlock_OPIN_84),
    .OPIN_85(logicBlock_OPIN_85),
    .OPIN_86(logicBlock_OPIN_86),
    .OPIN_87(logicBlock_OPIN_87),
    .OPIN_88(logicBlock_OPIN_88),
    .clock(logicBlock_clock),
    .reset(logicBlock_reset),
    .configBits(logicBlock_configBits),
    .loopBreak(logicBlock_loopBreak),
    .gndLBouts(logicBlock_gndLBouts)
  );
  ScanConf_Tile_7_1_clbmultile configBlock ( // @[TileFull.scala 66:31]
    .clock(configBlock_clock),
    .ioBundle_confOut(configBlock_ioBundle_confOut),
    .ioBundle_scan_in(configBlock_ioBundle_scan_in),
    .ioBundle_scan_en(configBlock_ioBundle_scan_en),
    .ioBundle_scan_out(configBlock_ioBundle_scan_out)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN0_N14762 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN0_N14762_io_in),
    .io_config(CBMux_IPIN0_N14762_io_config),
    .io_out(CBMux_IPIN0_N14762_io_out),
    .io_loopBreak(CBMux_IPIN0_N14762_io_loopBreak),
    .io_cnstClk(CBMux_IPIN0_N14762_io_cnstClk),
    .io_arst(CBMux_IPIN0_N14762_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN1_N14763 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN1_N14763_io_in),
    .io_config(CBMux_IPIN1_N14763_io_config),
    .io_out(CBMux_IPIN1_N14763_io_out),
    .io_loopBreak(CBMux_IPIN1_N14763_io_loopBreak),
    .io_cnstClk(CBMux_IPIN1_N14763_io_cnstClk),
    .io_arst(CBMux_IPIN1_N14763_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN2_N14764 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN2_N14764_io_in),
    .io_config(CBMux_IPIN2_N14764_io_config),
    .io_out(CBMux_IPIN2_N14764_io_out),
    .io_loopBreak(CBMux_IPIN2_N14764_io_loopBreak),
    .io_cnstClk(CBMux_IPIN2_N14764_io_cnstClk),
    .io_arst(CBMux_IPIN2_N14764_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN3_N14765 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN3_N14765_io_in),
    .io_config(CBMux_IPIN3_N14765_io_config),
    .io_out(CBMux_IPIN3_N14765_io_out),
    .io_loopBreak(CBMux_IPIN3_N14765_io_loopBreak),
    .io_cnstClk(CBMux_IPIN3_N14765_io_cnstClk),
    .io_arst(CBMux_IPIN3_N14765_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN4_N14766 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN4_N14766_io_in),
    .io_config(CBMux_IPIN4_N14766_io_config),
    .io_out(CBMux_IPIN4_N14766_io_out),
    .io_loopBreak(CBMux_IPIN4_N14766_io_loopBreak),
    .io_cnstClk(CBMux_IPIN4_N14766_io_cnstClk),
    .io_arst(CBMux_IPIN4_N14766_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN5_N14767 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN5_N14767_io_in),
    .io_config(CBMux_IPIN5_N14767_io_config),
    .io_out(CBMux_IPIN5_N14767_io_out),
    .io_loopBreak(CBMux_IPIN5_N14767_io_loopBreak),
    .io_cnstClk(CBMux_IPIN5_N14767_io_cnstClk),
    .io_arst(CBMux_IPIN5_N14767_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN6_N14768 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN6_N14768_io_in),
    .io_config(CBMux_IPIN6_N14768_io_config),
    .io_out(CBMux_IPIN6_N14768_io_out),
    .io_loopBreak(CBMux_IPIN6_N14768_io_loopBreak),
    .io_cnstClk(CBMux_IPIN6_N14768_io_cnstClk),
    .io_arst(CBMux_IPIN6_N14768_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN7_N14769 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN7_N14769_io_in),
    .io_config(CBMux_IPIN7_N14769_io_config),
    .io_out(CBMux_IPIN7_N14769_io_out),
    .io_loopBreak(CBMux_IPIN7_N14769_io_loopBreak),
    .io_cnstClk(CBMux_IPIN7_N14769_io_cnstClk),
    .io_arst(CBMux_IPIN7_N14769_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN8_N14770 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN8_N14770_io_in),
    .io_config(CBMux_IPIN8_N14770_io_config),
    .io_out(CBMux_IPIN8_N14770_io_out),
    .io_loopBreak(CBMux_IPIN8_N14770_io_loopBreak),
    .io_cnstClk(CBMux_IPIN8_N14770_io_cnstClk),
    .io_arst(CBMux_IPIN8_N14770_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN9_N14771 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN9_N14771_io_in),
    .io_config(CBMux_IPIN9_N14771_io_config),
    .io_out(CBMux_IPIN9_N14771_io_out),
    .io_loopBreak(CBMux_IPIN9_N14771_io_loopBreak),
    .io_cnstClk(CBMux_IPIN9_N14771_io_cnstClk),
    .io_arst(CBMux_IPIN9_N14771_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN10_N14772 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN10_N14772_io_in),
    .io_config(CBMux_IPIN10_N14772_io_config),
    .io_out(CBMux_IPIN10_N14772_io_out),
    .io_loopBreak(CBMux_IPIN10_N14772_io_loopBreak),
    .io_cnstClk(CBMux_IPIN10_N14772_io_cnstClk),
    .io_arst(CBMux_IPIN10_N14772_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN11_N14773 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN11_N14773_io_in),
    .io_config(CBMux_IPIN11_N14773_io_config),
    .io_out(CBMux_IPIN11_N14773_io_out),
    .io_loopBreak(CBMux_IPIN11_N14773_io_loopBreak),
    .io_cnstClk(CBMux_IPIN11_N14773_io_cnstClk),
    .io_arst(CBMux_IPIN11_N14773_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN12_N14774 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN12_N14774_io_in),
    .io_config(CBMux_IPIN12_N14774_io_config),
    .io_out(CBMux_IPIN12_N14774_io_out),
    .io_loopBreak(CBMux_IPIN12_N14774_io_loopBreak),
    .io_cnstClk(CBMux_IPIN12_N14774_io_cnstClk),
    .io_arst(CBMux_IPIN12_N14774_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN13_N14775 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN13_N14775_io_in),
    .io_config(CBMux_IPIN13_N14775_io_config),
    .io_out(CBMux_IPIN13_N14775_io_out),
    .io_loopBreak(CBMux_IPIN13_N14775_io_loopBreak),
    .io_cnstClk(CBMux_IPIN13_N14775_io_cnstClk),
    .io_arst(CBMux_IPIN13_N14775_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN14_N14776 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN14_N14776_io_in),
    .io_config(CBMux_IPIN14_N14776_io_config),
    .io_out(CBMux_IPIN14_N14776_io_out),
    .io_loopBreak(CBMux_IPIN14_N14776_io_loopBreak),
    .io_cnstClk(CBMux_IPIN14_N14776_io_cnstClk),
    .io_arst(CBMux_IPIN14_N14776_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN15_N14777 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN15_N14777_io_in),
    .io_config(CBMux_IPIN15_N14777_io_config),
    .io_out(CBMux_IPIN15_N14777_io_out),
    .io_loopBreak(CBMux_IPIN15_N14777_io_loopBreak),
    .io_cnstClk(CBMux_IPIN15_N14777_io_cnstClk),
    .io_arst(CBMux_IPIN15_N14777_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN16_N14778 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN16_N14778_io_in),
    .io_config(CBMux_IPIN16_N14778_io_config),
    .io_out(CBMux_IPIN16_N14778_io_out),
    .io_loopBreak(CBMux_IPIN16_N14778_io_loopBreak),
    .io_cnstClk(CBMux_IPIN16_N14778_io_cnstClk),
    .io_arst(CBMux_IPIN16_N14778_io_arst)
  );
  MuxNInput_28_SCAOptCB CBMux_IPIN17_N14779 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN17_N14779_io_in),
    .io_config(CBMux_IPIN17_N14779_io_config),
    .io_out(CBMux_IPIN17_N14779_io_out),
    .io_loopBreak(CBMux_IPIN17_N14779_io_loopBreak),
    .io_cnstClk(CBMux_IPIN17_N14779_io_cnstClk),
    .io_arst(CBMux_IPIN17_N14779_io_arst)
  );
  MuxNInput_24_SCAOptCB CBMux_IPIN18_N14780 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN18_N14780_io_in),
    .io_config(CBMux_IPIN18_N14780_io_config),
    .io_out(CBMux_IPIN18_N14780_io_out),
    .io_loopBreak(CBMux_IPIN18_N14780_io_loopBreak),
    .io_cnstClk(CBMux_IPIN18_N14780_io_cnstClk),
    .io_arst(CBMux_IPIN18_N14780_io_arst)
  );
  MuxNInput_24_SCAOptCB CBMux_IPIN19_N14781 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN19_N14781_io_in),
    .io_config(CBMux_IPIN19_N14781_io_config),
    .io_out(CBMux_IPIN19_N14781_io_out),
    .io_loopBreak(CBMux_IPIN19_N14781_io_loopBreak),
    .io_cnstClk(CBMux_IPIN19_N14781_io_cnstClk),
    .io_arst(CBMux_IPIN19_N14781_io_arst)
  );
  MuxNInput_22_SCAOptCB CBMux_IPIN20_N14782 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN20_N14782_io_in),
    .io_config(CBMux_IPIN20_N14782_io_config),
    .io_out(CBMux_IPIN20_N14782_io_out),
    .io_loopBreak(CBMux_IPIN20_N14782_io_loopBreak),
    .io_cnstClk(CBMux_IPIN20_N14782_io_cnstClk),
    .io_arst(CBMux_IPIN20_N14782_io_arst)
  );
  MuxNInput_26_SCAOptCB CBMux_IPIN21_N14783 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN21_N14783_io_in),
    .io_config(CBMux_IPIN21_N14783_io_config),
    .io_out(CBMux_IPIN21_N14783_io_out),
    .io_loopBreak(CBMux_IPIN21_N14783_io_loopBreak),
    .io_cnstClk(CBMux_IPIN21_N14783_io_cnstClk),
    .io_arst(CBMux_IPIN21_N14783_io_arst)
  );
  MuxNInput_26_SCAOptCB CBMux_IPIN22_N14784 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN22_N14784_io_in),
    .io_config(CBMux_IPIN22_N14784_io_config),
    .io_out(CBMux_IPIN22_N14784_io_out),
    .io_loopBreak(CBMux_IPIN22_N14784_io_loopBreak),
    .io_cnstClk(CBMux_IPIN22_N14784_io_cnstClk),
    .io_arst(CBMux_IPIN22_N14784_io_arst)
  );
  MuxNInput_22_SCAOptCB CBMux_IPIN23_N14785 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN23_N14785_io_in),
    .io_config(CBMux_IPIN23_N14785_io_config),
    .io_out(CBMux_IPIN23_N14785_io_out),
    .io_loopBreak(CBMux_IPIN23_N14785_io_loopBreak),
    .io_cnstClk(CBMux_IPIN23_N14785_io_cnstClk),
    .io_arst(CBMux_IPIN23_N14785_io_arst)
  );
  MuxNInput_22_SCAOptCB CBMux_IPIN24_N14786 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN24_N14786_io_in),
    .io_config(CBMux_IPIN24_N14786_io_config),
    .io_out(CBMux_IPIN24_N14786_io_out),
    .io_loopBreak(CBMux_IPIN24_N14786_io_loopBreak),
    .io_cnstClk(CBMux_IPIN24_N14786_io_cnstClk),
    .io_arst(CBMux_IPIN24_N14786_io_arst)
  );
  MuxNInput_22_SCAOptCB CBMux_IPIN25_N14787 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN25_N14787_io_in),
    .io_config(CBMux_IPIN25_N14787_io_config),
    .io_out(CBMux_IPIN25_N14787_io_out),
    .io_loopBreak(CBMux_IPIN25_N14787_io_loopBreak),
    .io_cnstClk(CBMux_IPIN25_N14787_io_cnstClk),
    .io_arst(CBMux_IPIN25_N14787_io_arst)
  );
  MuxNInput_26_SCAOptCB CBMux_IPIN26_N14788 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN26_N14788_io_in),
    .io_config(CBMux_IPIN26_N14788_io_config),
    .io_out(CBMux_IPIN26_N14788_io_out),
    .io_loopBreak(CBMux_IPIN26_N14788_io_loopBreak),
    .io_cnstClk(CBMux_IPIN26_N14788_io_cnstClk),
    .io_arst(CBMux_IPIN26_N14788_io_arst)
  );
  MuxNInput_26_SCAOptCB CBMux_IPIN27_N14789 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN27_N14789_io_in),
    .io_config(CBMux_IPIN27_N14789_io_config),
    .io_out(CBMux_IPIN27_N14789_io_out),
    .io_loopBreak(CBMux_IPIN27_N14789_io_loopBreak),
    .io_cnstClk(CBMux_IPIN27_N14789_io_cnstClk),
    .io_arst(CBMux_IPIN27_N14789_io_arst)
  );
  MuxNInput_26_SCAOptCB CBMux_IPIN28_N14790 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN28_N14790_io_in),
    .io_config(CBMux_IPIN28_N14790_io_config),
    .io_out(CBMux_IPIN28_N14790_io_out),
    .io_loopBreak(CBMux_IPIN28_N14790_io_loopBreak),
    .io_cnstClk(CBMux_IPIN28_N14790_io_cnstClk),
    .io_arst(CBMux_IPIN28_N14790_io_arst)
  );
  MuxNInput_22_SCAOptCB CBMux_IPIN29_N14791 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN29_N14791_io_in),
    .io_config(CBMux_IPIN29_N14791_io_config),
    .io_out(CBMux_IPIN29_N14791_io_out),
    .io_loopBreak(CBMux_IPIN29_N14791_io_loopBreak),
    .io_cnstClk(CBMux_IPIN29_N14791_io_cnstClk),
    .io_arst(CBMux_IPIN29_N14791_io_arst)
  );
  MuxNInput_22_SCAOptCB CBMux_IPIN30_N14792 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN30_N14792_io_in),
    .io_config(CBMux_IPIN30_N14792_io_config),
    .io_out(CBMux_IPIN30_N14792_io_out),
    .io_loopBreak(CBMux_IPIN30_N14792_io_loopBreak),
    .io_cnstClk(CBMux_IPIN30_N14792_io_cnstClk),
    .io_arst(CBMux_IPIN30_N14792_io_arst)
  );
  MuxNInput_26_SCAOptCB CBMux_IPIN31_N14793 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN31_N14793_io_in),
    .io_config(CBMux_IPIN31_N14793_io_config),
    .io_out(CBMux_IPIN31_N14793_io_out),
    .io_loopBreak(CBMux_IPIN31_N14793_io_loopBreak),
    .io_cnstClk(CBMux_IPIN31_N14793_io_cnstClk),
    .io_arst(CBMux_IPIN31_N14793_io_arst)
  );
  MuxNInput_26_SCAOptCB CBMux_IPIN32_N14794 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN32_N14794_io_in),
    .io_config(CBMux_IPIN32_N14794_io_config),
    .io_out(CBMux_IPIN32_N14794_io_out),
    .io_loopBreak(CBMux_IPIN32_N14794_io_loopBreak),
    .io_cnstClk(CBMux_IPIN32_N14794_io_cnstClk),
    .io_arst(CBMux_IPIN32_N14794_io_arst)
  );
  MuxNInput_26_SCAOptCB CBMux_IPIN33_N14795 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN33_N14795_io_in),
    .io_config(CBMux_IPIN33_N14795_io_config),
    .io_out(CBMux_IPIN33_N14795_io_out),
    .io_loopBreak(CBMux_IPIN33_N14795_io_loopBreak),
    .io_cnstClk(CBMux_IPIN33_N14795_io_cnstClk),
    .io_arst(CBMux_IPIN33_N14795_io_arst)
  );
  MuxNInput_22_SCAOptCB CBMux_IPIN34_N14796 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN34_N14796_io_in),
    .io_config(CBMux_IPIN34_N14796_io_config),
    .io_out(CBMux_IPIN34_N14796_io_out),
    .io_loopBreak(CBMux_IPIN34_N14796_io_loopBreak),
    .io_cnstClk(CBMux_IPIN34_N14796_io_cnstClk),
    .io_arst(CBMux_IPIN34_N14796_io_arst)
  );
  MuxNInput_22_SCAOptCB CBMux_IPIN35_N14797 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN35_N14797_io_in),
    .io_config(CBMux_IPIN35_N14797_io_config),
    .io_out(CBMux_IPIN35_N14797_io_out),
    .io_loopBreak(CBMux_IPIN35_N14797_io_loopBreak),
    .io_cnstClk(CBMux_IPIN35_N14797_io_cnstClk),
    .io_arst(CBMux_IPIN35_N14797_io_arst)
  );
  MuxNInput_22_SCAOptCB CBMux_IPIN36_N14798 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN36_N14798_io_in),
    .io_config(CBMux_IPIN36_N14798_io_config),
    .io_out(CBMux_IPIN36_N14798_io_out),
    .io_loopBreak(CBMux_IPIN36_N14798_io_loopBreak),
    .io_cnstClk(CBMux_IPIN36_N14798_io_cnstClk),
    .io_arst(CBMux_IPIN36_N14798_io_arst)
  );
  MuxNInput_26_SCAOptCB CBMux_IPIN37_N14799 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN37_N14799_io_in),
    .io_config(CBMux_IPIN37_N14799_io_config),
    .io_out(CBMux_IPIN37_N14799_io_out),
    .io_loopBreak(CBMux_IPIN37_N14799_io_loopBreak),
    .io_cnstClk(CBMux_IPIN37_N14799_io_cnstClk),
    .io_arst(CBMux_IPIN37_N14799_io_arst)
  );
  MuxNInput_26_SCAOptCB CBMux_IPIN38_N14800 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN38_N14800_io_in),
    .io_config(CBMux_IPIN38_N14800_io_config),
    .io_out(CBMux_IPIN38_N14800_io_out),
    .io_loopBreak(CBMux_IPIN38_N14800_io_loopBreak),
    .io_cnstClk(CBMux_IPIN38_N14800_io_cnstClk),
    .io_arst(CBMux_IPIN38_N14800_io_arst)
  );
  MuxNInput_22_SCAOptCB CBMux_IPIN39_N14801 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN39_N14801_io_in),
    .io_config(CBMux_IPIN39_N14801_io_config),
    .io_out(CBMux_IPIN39_N14801_io_out),
    .io_loopBreak(CBMux_IPIN39_N14801_io_loopBreak),
    .io_cnstClk(CBMux_IPIN39_N14801_io_cnstClk),
    .io_arst(CBMux_IPIN39_N14801_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN40_N14802 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN40_N14802_io_in),
    .io_config(CBMux_IPIN40_N14802_io_config),
    .io_out(CBMux_IPIN40_N14802_io_out),
    .io_loopBreak(CBMux_IPIN40_N14802_io_loopBreak),
    .io_cnstClk(CBMux_IPIN40_N14802_io_cnstClk),
    .io_arst(CBMux_IPIN40_N14802_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN41_N14803 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN41_N14803_io_in),
    .io_config(CBMux_IPIN41_N14803_io_config),
    .io_out(CBMux_IPIN41_N14803_io_out),
    .io_loopBreak(CBMux_IPIN41_N14803_io_loopBreak),
    .io_cnstClk(CBMux_IPIN41_N14803_io_cnstClk),
    .io_arst(CBMux_IPIN41_N14803_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN42_N14804 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN42_N14804_io_in),
    .io_config(CBMux_IPIN42_N14804_io_config),
    .io_out(CBMux_IPIN42_N14804_io_out),
    .io_loopBreak(CBMux_IPIN42_N14804_io_loopBreak),
    .io_cnstClk(CBMux_IPIN42_N14804_io_cnstClk),
    .io_arst(CBMux_IPIN42_N14804_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN43_N14805 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN43_N14805_io_in),
    .io_config(CBMux_IPIN43_N14805_io_config),
    .io_out(CBMux_IPIN43_N14805_io_out),
    .io_loopBreak(CBMux_IPIN43_N14805_io_loopBreak),
    .io_cnstClk(CBMux_IPIN43_N14805_io_cnstClk),
    .io_arst(CBMux_IPIN43_N14805_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN44_N14806 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN44_N14806_io_in),
    .io_config(CBMux_IPIN44_N14806_io_config),
    .io_out(CBMux_IPIN44_N14806_io_out),
    .io_loopBreak(CBMux_IPIN44_N14806_io_loopBreak),
    .io_cnstClk(CBMux_IPIN44_N14806_io_cnstClk),
    .io_arst(CBMux_IPIN44_N14806_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN45_N14807 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN45_N14807_io_in),
    .io_config(CBMux_IPIN45_N14807_io_config),
    .io_out(CBMux_IPIN45_N14807_io_out),
    .io_loopBreak(CBMux_IPIN45_N14807_io_loopBreak),
    .io_cnstClk(CBMux_IPIN45_N14807_io_cnstClk),
    .io_arst(CBMux_IPIN45_N14807_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN46_N14808 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN46_N14808_io_in),
    .io_config(CBMux_IPIN46_N14808_io_config),
    .io_out(CBMux_IPIN46_N14808_io_out),
    .io_loopBreak(CBMux_IPIN46_N14808_io_loopBreak),
    .io_cnstClk(CBMux_IPIN46_N14808_io_cnstClk),
    .io_arst(CBMux_IPIN46_N14808_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN47_N14809 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN47_N14809_io_in),
    .io_config(CBMux_IPIN47_N14809_io_config),
    .io_out(CBMux_IPIN47_N14809_io_out),
    .io_loopBreak(CBMux_IPIN47_N14809_io_loopBreak),
    .io_cnstClk(CBMux_IPIN47_N14809_io_cnstClk),
    .io_arst(CBMux_IPIN47_N14809_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN48_N14810 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN48_N14810_io_in),
    .io_config(CBMux_IPIN48_N14810_io_config),
    .io_out(CBMux_IPIN48_N14810_io_out),
    .io_loopBreak(CBMux_IPIN48_N14810_io_loopBreak),
    .io_cnstClk(CBMux_IPIN48_N14810_io_cnstClk),
    .io_arst(CBMux_IPIN48_N14810_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN49_N14811 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN49_N14811_io_in),
    .io_config(CBMux_IPIN49_N14811_io_config),
    .io_out(CBMux_IPIN49_N14811_io_out),
    .io_loopBreak(CBMux_IPIN49_N14811_io_loopBreak),
    .io_cnstClk(CBMux_IPIN49_N14811_io_cnstClk),
    .io_arst(CBMux_IPIN49_N14811_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN50_N14812 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN50_N14812_io_in),
    .io_config(CBMux_IPIN50_N14812_io_config),
    .io_out(CBMux_IPIN50_N14812_io_out),
    .io_loopBreak(CBMux_IPIN50_N14812_io_loopBreak),
    .io_cnstClk(CBMux_IPIN50_N14812_io_cnstClk),
    .io_arst(CBMux_IPIN50_N14812_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN51_N14813 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN51_N14813_io_in),
    .io_config(CBMux_IPIN51_N14813_io_config),
    .io_out(CBMux_IPIN51_N14813_io_out),
    .io_loopBreak(CBMux_IPIN51_N14813_io_loopBreak),
    .io_cnstClk(CBMux_IPIN51_N14813_io_cnstClk),
    .io_arst(CBMux_IPIN51_N14813_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN52_N14814 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN52_N14814_io_in),
    .io_config(CBMux_IPIN52_N14814_io_config),
    .io_out(CBMux_IPIN52_N14814_io_out),
    .io_loopBreak(CBMux_IPIN52_N14814_io_loopBreak),
    .io_cnstClk(CBMux_IPIN52_N14814_io_cnstClk),
    .io_arst(CBMux_IPIN52_N14814_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN53_N14815 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN53_N14815_io_in),
    .io_config(CBMux_IPIN53_N14815_io_config),
    .io_out(CBMux_IPIN53_N14815_io_out),
    .io_loopBreak(CBMux_IPIN53_N14815_io_loopBreak),
    .io_cnstClk(CBMux_IPIN53_N14815_io_cnstClk),
    .io_arst(CBMux_IPIN53_N14815_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN54_N14816 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN54_N14816_io_in),
    .io_config(CBMux_IPIN54_N14816_io_config),
    .io_out(CBMux_IPIN54_N14816_io_out),
    .io_loopBreak(CBMux_IPIN54_N14816_io_loopBreak),
    .io_cnstClk(CBMux_IPIN54_N14816_io_cnstClk),
    .io_arst(CBMux_IPIN54_N14816_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN55_N14817 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN55_N14817_io_in),
    .io_config(CBMux_IPIN55_N14817_io_config),
    .io_out(CBMux_IPIN55_N14817_io_out),
    .io_loopBreak(CBMux_IPIN55_N14817_io_loopBreak),
    .io_cnstClk(CBMux_IPIN55_N14817_io_cnstClk),
    .io_arst(CBMux_IPIN55_N14817_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN56_N14818 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN56_N14818_io_in),
    .io_config(CBMux_IPIN56_N14818_io_config),
    .io_out(CBMux_IPIN56_N14818_io_out),
    .io_loopBreak(CBMux_IPIN56_N14818_io_loopBreak),
    .io_cnstClk(CBMux_IPIN56_N14818_io_cnstClk),
    .io_arst(CBMux_IPIN56_N14818_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN57_N14819 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN57_N14819_io_in),
    .io_config(CBMux_IPIN57_N14819_io_config),
    .io_out(CBMux_IPIN57_N14819_io_out),
    .io_loopBreak(CBMux_IPIN57_N14819_io_loopBreak),
    .io_cnstClk(CBMux_IPIN57_N14819_io_cnstClk),
    .io_arst(CBMux_IPIN57_N14819_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN58_N14820 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN58_N14820_io_in),
    .io_config(CBMux_IPIN58_N14820_io_config),
    .io_out(CBMux_IPIN58_N14820_io_out),
    .io_loopBreak(CBMux_IPIN58_N14820_io_loopBreak),
    .io_cnstClk(CBMux_IPIN58_N14820_io_cnstClk),
    .io_arst(CBMux_IPIN58_N14820_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN59_N14821 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN59_N14821_io_in),
    .io_config(CBMux_IPIN59_N14821_io_config),
    .io_out(CBMux_IPIN59_N14821_io_out),
    .io_loopBreak(CBMux_IPIN59_N14821_io_loopBreak),
    .io_cnstClk(CBMux_IPIN59_N14821_io_cnstClk),
    .io_arst(CBMux_IPIN59_N14821_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN60_N14822 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN60_N14822_io_in),
    .io_config(CBMux_IPIN60_N14822_io_config),
    .io_out(CBMux_IPIN60_N14822_io_out),
    .io_loopBreak(CBMux_IPIN60_N14822_io_loopBreak),
    .io_cnstClk(CBMux_IPIN60_N14822_io_cnstClk),
    .io_arst(CBMux_IPIN60_N14822_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN61_N14823 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN61_N14823_io_in),
    .io_config(CBMux_IPIN61_N14823_io_config),
    .io_out(CBMux_IPIN61_N14823_io_out),
    .io_loopBreak(CBMux_IPIN61_N14823_io_loopBreak),
    .io_cnstClk(CBMux_IPIN61_N14823_io_cnstClk),
    .io_arst(CBMux_IPIN61_N14823_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN62_N14824 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN62_N14824_io_in),
    .io_config(CBMux_IPIN62_N14824_io_config),
    .io_out(CBMux_IPIN62_N14824_io_out),
    .io_loopBreak(CBMux_IPIN62_N14824_io_loopBreak),
    .io_cnstClk(CBMux_IPIN62_N14824_io_cnstClk),
    .io_arst(CBMux_IPIN62_N14824_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN63_N14825 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN63_N14825_io_in),
    .io_config(CBMux_IPIN63_N14825_io_config),
    .io_out(CBMux_IPIN63_N14825_io_out),
    .io_loopBreak(CBMux_IPIN63_N14825_io_loopBreak),
    .io_cnstClk(CBMux_IPIN63_N14825_io_cnstClk),
    .io_arst(CBMux_IPIN63_N14825_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN64_N14826 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN64_N14826_io_in),
    .io_config(CBMux_IPIN64_N14826_io_config),
    .io_out(CBMux_IPIN64_N14826_io_out),
    .io_loopBreak(CBMux_IPIN64_N14826_io_loopBreak),
    .io_cnstClk(CBMux_IPIN64_N14826_io_cnstClk),
    .io_arst(CBMux_IPIN64_N14826_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN65_N14827 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN65_N14827_io_in),
    .io_config(CBMux_IPIN65_N14827_io_config),
    .io_out(CBMux_IPIN65_N14827_io_out),
    .io_loopBreak(CBMux_IPIN65_N14827_io_loopBreak),
    .io_cnstClk(CBMux_IPIN65_N14827_io_cnstClk),
    .io_arst(CBMux_IPIN65_N14827_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN66_N14828 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN66_N14828_io_in),
    .io_config(CBMux_IPIN66_N14828_io_config),
    .io_out(CBMux_IPIN66_N14828_io_out),
    .io_loopBreak(CBMux_IPIN66_N14828_io_loopBreak),
    .io_cnstClk(CBMux_IPIN66_N14828_io_cnstClk),
    .io_arst(CBMux_IPIN66_N14828_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN67_N14829 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN67_N14829_io_in),
    .io_config(CBMux_IPIN67_N14829_io_config),
    .io_out(CBMux_IPIN67_N14829_io_out),
    .io_loopBreak(CBMux_IPIN67_N14829_io_loopBreak),
    .io_cnstClk(CBMux_IPIN67_N14829_io_cnstClk),
    .io_arst(CBMux_IPIN67_N14829_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN68_N14830 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN68_N14830_io_in),
    .io_config(CBMux_IPIN68_N14830_io_config),
    .io_out(CBMux_IPIN68_N14830_io_out),
    .io_loopBreak(CBMux_IPIN68_N14830_io_loopBreak),
    .io_cnstClk(CBMux_IPIN68_N14830_io_cnstClk),
    .io_arst(CBMux_IPIN68_N14830_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN69_N14831 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN69_N14831_io_in),
    .io_config(CBMux_IPIN69_N14831_io_config),
    .io_out(CBMux_IPIN69_N14831_io_out),
    .io_loopBreak(CBMux_IPIN69_N14831_io_loopBreak),
    .io_cnstClk(CBMux_IPIN69_N14831_io_cnstClk),
    .io_arst(CBMux_IPIN69_N14831_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN70_N14832 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN70_N14832_io_in),
    .io_config(CBMux_IPIN70_N14832_io_config),
    .io_out(CBMux_IPIN70_N14832_io_out),
    .io_loopBreak(CBMux_IPIN70_N14832_io_loopBreak),
    .io_cnstClk(CBMux_IPIN70_N14832_io_cnstClk),
    .io_arst(CBMux_IPIN70_N14832_io_arst)
  );
  MuxNInput_1_SCAOptCB CBMux_IPIN71_N14833 ( // @[TileFull.scala 102:29]
    .io_in(CBMux_IPIN71_N14833_io_in),
    .io_config(CBMux_IPIN71_N14833_io_config),
    .io_out(CBMux_IPIN71_N14833_io_out),
    .io_loopBreak(CBMux_IPIN71_N14833_io_loopBreak),
    .io_cnstClk(CBMux_IPIN71_N14833_io_cnstClk),
    .io_arst(CBMux_IPIN71_N14833_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C1_N23683_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C1_N23683_O_3_C_6_io_in),
    .io_config(SBMux_C1_N23683_O_3_C_6_io_config),
    .io_out(SBMux_C1_N23683_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C1_N23683_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C1_N23683_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C1_N23683_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C1_N23683_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C7_SCAOptSB SBMux_C9_N23685_O_3_C_7 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C9_N23685_O_3_C_7_io_in),
    .io_config(SBMux_C9_N23685_O_3_C_7_io_config),
    .io_out(SBMux_C9_N23685_O_3_C_7_io_out),
    .io_loopBreak(SBMux_C9_N23685_O_3_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C9_N23685_O_3_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C9_N23685_O_3_C_7_io_cnstClk),
    .io_arst(SBMux_C9_N23685_O_3_C_7_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C17_N23687_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C17_N23687_O_3_C_6_io_in),
    .io_config(SBMux_C17_N23687_O_3_C_6_io_config),
    .io_out(SBMux_C17_N23687_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C17_N23687_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C17_N23687_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C17_N23687_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C17_N23687_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C25_N23689_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C25_N23689_O_3_C_6_io_in),
    .io_config(SBMux_C25_N23689_O_3_C_6_io_config),
    .io_out(SBMux_C25_N23689_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C25_N23689_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C25_N23689_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C25_N23689_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C25_N23689_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C7_SCAOptSB SBMux_C33_N23691_O_3_C_7 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C33_N23691_O_3_C_7_io_in),
    .io_config(SBMux_C33_N23691_O_3_C_7_io_config),
    .io_out(SBMux_C33_N23691_O_3_C_7_io_out),
    .io_loopBreak(SBMux_C33_N23691_O_3_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C33_N23691_O_3_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C33_N23691_O_3_C_7_io_cnstClk),
    .io_arst(SBMux_C33_N23691_O_3_C_7_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C41_N23693_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C41_N23693_O_3_C_6_io_in),
    .io_config(SBMux_C41_N23693_O_3_C_6_io_config),
    .io_out(SBMux_C41_N23693_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C41_N23693_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C41_N23693_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C41_N23693_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C41_N23693_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C49_N23695_O_3_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C49_N23695_O_3_C_5_io_in),
    .io_config(SBMux_C49_N23695_O_3_C_5_io_config),
    .io_out(SBMux_C49_N23695_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C49_N23695_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C49_N23695_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C49_N23695_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C49_N23695_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C57_N23697_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C57_N23697_O_3_C_6_io_in),
    .io_config(SBMux_C57_N23697_O_3_C_6_io_config),
    .io_out(SBMux_C57_N23697_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C57_N23697_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C57_N23697_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C57_N23697_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C57_N23697_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C65_N23699_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C65_N23699_O_3_C_6_io_in),
    .io_config(SBMux_C65_N23699_O_3_C_6_io_config),
    .io_out(SBMux_C65_N23699_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C65_N23699_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C65_N23699_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C65_N23699_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C65_N23699_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C73_N23701_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C73_N23701_O_3_C_6_io_in),
    .io_config(SBMux_C73_N23701_O_3_C_6_io_config),
    .io_out(SBMux_C73_N23701_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C73_N23701_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C73_N23701_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C73_N23701_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C73_N23701_O_3_C_6_io_arst)
  );
  MuxNInput_O2_C5_SCAOptSB SBMux_C81_N23703_O_2_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C81_N23703_O_2_C_5_io_in),
    .io_config(SBMux_C81_N23703_O_2_C_5_io_config),
    .io_out(SBMux_C81_N23703_O_2_C_5_io_out),
    .io_loopBreak(SBMux_C81_N23703_O_2_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C81_N23703_O_2_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C81_N23703_O_2_C_5_io_cnstClk),
    .io_arst(SBMux_C81_N23703_O_2_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C89_N23705_O_3_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C89_N23705_O_3_C_5_io_in),
    .io_config(SBMux_C89_N23705_O_3_C_5_io_config),
    .io_out(SBMux_C89_N23705_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C89_N23705_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C89_N23705_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C89_N23705_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C89_N23705_O_3_C_5_io_arst)
  );
  MuxNInput_O2_C5_SCAOptSB SBMux_C97_N23707_O_2_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C97_N23707_O_2_C_5_io_in),
    .io_config(SBMux_C97_N23707_O_2_C_5_io_config),
    .io_out(SBMux_C97_N23707_O_2_C_5_io_out),
    .io_loopBreak(SBMux_C97_N23707_O_2_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C97_N23707_O_2_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C97_N23707_O_2_C_5_io_cnstClk),
    .io_arst(SBMux_C97_N23707_O_2_C_5_io_arst)
  );
  MuxNInput_O0_C1_SCAOptSB SBMux_C101_N23767_O_0_C_1 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C101_N23767_O_0_C_1_io_in),
    .io_config(SBMux_C101_N23767_O_0_C_1_io_config),
    .io_out(SBMux_C101_N23767_O_0_C_1_io_out),
    .io_loopBreak(SBMux_C101_N23767_O_0_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C101_N23767_O_0_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C101_N23767_O_0_C_1_io_cnstClk),
    .io_arst(SBMux_C101_N23767_O_0_C_1_io_arst)
  );
  MuxNInput_O0_C1_SCAOptSB SBMux_C105_N23769_O_0_C_1 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C105_N23769_O_0_C_1_io_in),
    .io_config(SBMux_C105_N23769_O_0_C_1_io_config),
    .io_out(SBMux_C105_N23769_O_0_C_1_io_out),
    .io_loopBreak(SBMux_C105_N23769_O_0_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C105_N23769_O_0_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C105_N23769_O_0_C_1_io_cnstClk),
    .io_arst(SBMux_C105_N23769_O_0_C_1_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C0_N23798_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C0_N23798_O_3_C_6_io_in),
    .io_config(SBMux_C0_N23798_O_3_C_6_io_config),
    .io_out(SBMux_C0_N23798_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C0_N23798_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C0_N23798_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C0_N23798_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C0_N23798_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C8_N23800_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C8_N23800_O_3_C_6_io_in),
    .io_config(SBMux_C8_N23800_O_3_C_6_io_config),
    .io_out(SBMux_C8_N23800_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C8_N23800_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C8_N23800_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C8_N23800_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C8_N23800_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C16_N23802_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C16_N23802_O_3_C_6_io_in),
    .io_config(SBMux_C16_N23802_O_3_C_6_io_config),
    .io_out(SBMux_C16_N23802_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C16_N23802_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C16_N23802_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C16_N23802_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C16_N23802_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C7_SCAOptSB SBMux_C24_N23804_O_3_C_7 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C24_N23804_O_3_C_7_io_in),
    .io_config(SBMux_C24_N23804_O_3_C_7_io_config),
    .io_out(SBMux_C24_N23804_O_3_C_7_io_out),
    .io_loopBreak(SBMux_C24_N23804_O_3_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C24_N23804_O_3_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C24_N23804_O_3_C_7_io_cnstClk),
    .io_arst(SBMux_C24_N23804_O_3_C_7_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C32_N23806_O_3_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C32_N23806_O_3_C_5_io_in),
    .io_config(SBMux_C32_N23806_O_3_C_5_io_config),
    .io_out(SBMux_C32_N23806_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C32_N23806_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C32_N23806_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C32_N23806_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C32_N23806_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C40_N23808_O_3_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C40_N23808_O_3_C_5_io_in),
    .io_config(SBMux_C40_N23808_O_3_C_5_io_config),
    .io_out(SBMux_C40_N23808_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C40_N23808_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C40_N23808_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C40_N23808_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C40_N23808_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C48_N23810_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C48_N23810_O_3_C_6_io_in),
    .io_config(SBMux_C48_N23810_O_3_C_6_io_config),
    .io_out(SBMux_C48_N23810_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C48_N23810_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C48_N23810_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C48_N23810_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C48_N23810_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C56_N23812_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C56_N23812_O_3_C_6_io_in),
    .io_config(SBMux_C56_N23812_O_3_C_6_io_config),
    .io_out(SBMux_C56_N23812_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C56_N23812_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C56_N23812_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C56_N23812_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C56_N23812_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C64_N23814_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C64_N23814_O_3_C_6_io_in),
    .io_config(SBMux_C64_N23814_O_3_C_6_io_config),
    .io_out(SBMux_C64_N23814_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C64_N23814_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C64_N23814_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C64_N23814_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C64_N23814_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C7_SCAOptSB SBMux_C72_N23816_O_3_C_7 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C72_N23816_O_3_C_7_io_in),
    .io_config(SBMux_C72_N23816_O_3_C_7_io_config),
    .io_out(SBMux_C72_N23816_O_3_C_7_io_out),
    .io_loopBreak(SBMux_C72_N23816_O_3_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C72_N23816_O_3_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C72_N23816_O_3_C_7_io_cnstClk),
    .io_arst(SBMux_C72_N23816_O_3_C_7_io_arst)
  );
  MuxNInput_O2_C6_SCAOptSB SBMux_C80_N23818_O_2_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C80_N23818_O_2_C_6_io_in),
    .io_config(SBMux_C80_N23818_O_2_C_6_io_config),
    .io_out(SBMux_C80_N23818_O_2_C_6_io_out),
    .io_loopBreak(SBMux_C80_N23818_O_2_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C80_N23818_O_2_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C80_N23818_O_2_C_6_io_cnstClk),
    .io_arst(SBMux_C80_N23818_O_2_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C88_N23820_O_3_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C88_N23820_O_3_C_5_io_in),
    .io_config(SBMux_C88_N23820_O_3_C_5_io_config),
    .io_out(SBMux_C88_N23820_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C88_N23820_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C88_N23820_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C88_N23820_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C88_N23820_O_3_C_5_io_arst)
  );
  MuxNInput_O2_C5_SCAOptSB SBMux_C96_N23822_O_2_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C96_N23822_O_2_C_5_io_in),
    .io_config(SBMux_C96_N23822_O_2_C_5_io_config),
    .io_out(SBMux_C96_N23822_O_2_C_5_io_out),
    .io_loopBreak(SBMux_C96_N23822_O_2_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C96_N23822_O_2_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C96_N23822_O_2_C_5_io_cnstClk),
    .io_arst(SBMux_C96_N23822_O_2_C_5_io_arst)
  );
  MuxNInput_O0_C1_SCAOptSB SBMux_C100_N23824_O_0_C_1 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C100_N23824_O_0_C_1_io_in),
    .io_config(SBMux_C100_N23824_O_0_C_1_io_config),
    .io_out(SBMux_C100_N23824_O_0_C_1_io_out),
    .io_loopBreak(SBMux_C100_N23824_O_0_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C100_N23824_O_0_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C100_N23824_O_0_C_1_io_cnstClk),
    .io_arst(SBMux_C100_N23824_O_0_C_1_io_arst)
  );
  MuxNInput_O0_C1_SCAOptSB SBMux_C104_N23826_O_0_C_1 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C104_N23826_O_0_C_1_io_in),
    .io_config(SBMux_C104_N23826_O_0_C_1_io_config),
    .io_out(SBMux_C104_N23826_O_0_C_1_io_out),
    .io_loopBreak(SBMux_C104_N23826_O_0_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C104_N23826_O_0_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C104_N23826_O_0_C_1_io_cnstClk),
    .io_arst(SBMux_C104_N23826_O_0_C_1_io_arst)
  );
  MuxNInput_O4_C6_SCAOptSB SBMux_C1_N30079_O_4_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C1_N30079_O_4_C_6_io_in),
    .io_config(SBMux_C1_N30079_O_4_C_6_io_config),
    .io_out(SBMux_C1_N30079_O_4_C_6_io_out),
    .io_loopBreak(SBMux_C1_N30079_O_4_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C1_N30079_O_4_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C1_N30079_O_4_C_6_io_cnstClk),
    .io_arst(SBMux_C1_N30079_O_4_C_6_io_arst)
  );
  MuxNInput_O4_C7_SCAOptSB SBMux_C9_N30087_O_4_C_7 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C9_N30087_O_4_C_7_io_in),
    .io_config(SBMux_C9_N30087_O_4_C_7_io_config),
    .io_out(SBMux_C9_N30087_O_4_C_7_io_out),
    .io_loopBreak(SBMux_C9_N30087_O_4_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C9_N30087_O_4_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C9_N30087_O_4_C_7_io_cnstClk),
    .io_arst(SBMux_C9_N30087_O_4_C_7_io_arst)
  );
  MuxNInput_O3_C7_SCAOptSB SBMux_C17_N30095_O_3_C_7 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C17_N30095_O_3_C_7_io_in),
    .io_config(SBMux_C17_N30095_O_3_C_7_io_config),
    .io_out(SBMux_C17_N30095_O_3_C_7_io_out),
    .io_loopBreak(SBMux_C17_N30095_O_3_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C17_N30095_O_3_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C17_N30095_O_3_C_7_io_cnstClk),
    .io_arst(SBMux_C17_N30095_O_3_C_7_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C25_N30103_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C25_N30103_O_3_C_6_io_in),
    .io_config(SBMux_C25_N30103_O_3_C_6_io_config),
    .io_out(SBMux_C25_N30103_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C25_N30103_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C25_N30103_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C25_N30103_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C25_N30103_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C4_SCAOptSB SBMux_C33_N30111_O_3_C_4 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C33_N30111_O_3_C_4_io_in),
    .io_config(SBMux_C33_N30111_O_3_C_4_io_config),
    .io_out(SBMux_C33_N30111_O_3_C_4_io_out),
    .io_loopBreak(SBMux_C33_N30111_O_3_C_4_io_loopBreak),
    .io_ioGndBle(SBMux_C33_N30111_O_3_C_4_io_ioGndBle),
    .io_cnstClk(SBMux_C33_N30111_O_3_C_4_io_cnstClk),
    .io_arst(SBMux_C33_N30111_O_3_C_4_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C41_N30119_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C41_N30119_O_3_C_6_io_in),
    .io_config(SBMux_C41_N30119_O_3_C_6_io_config),
    .io_out(SBMux_C41_N30119_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C41_N30119_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C41_N30119_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C41_N30119_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C41_N30119_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C49_N30127_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C49_N30127_O_3_C_6_io_in),
    .io_config(SBMux_C49_N30127_O_3_C_6_io_config),
    .io_out(SBMux_C49_N30127_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C49_N30127_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C49_N30127_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C49_N30127_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C49_N30127_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C57_N30135_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C57_N30135_O_3_C_6_io_in),
    .io_config(SBMux_C57_N30135_O_3_C_6_io_config),
    .io_out(SBMux_C57_N30135_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C57_N30135_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C57_N30135_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C57_N30135_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C57_N30135_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C65_N30143_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C65_N30143_O_3_C_6_io_in),
    .io_config(SBMux_C65_N30143_O_3_C_6_io_config),
    .io_out(SBMux_C65_N30143_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C65_N30143_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C65_N30143_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C65_N30143_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C65_N30143_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C73_N30151_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C73_N30151_O_3_C_6_io_in),
    .io_config(SBMux_C73_N30151_O_3_C_6_io_config),
    .io_out(SBMux_C73_N30151_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C73_N30151_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C73_N30151_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C73_N30151_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C73_N30151_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C81_N30159_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C81_N30159_O_3_C_6_io_in),
    .io_config(SBMux_C81_N30159_O_3_C_6_io_config),
    .io_out(SBMux_C81_N30159_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C81_N30159_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C81_N30159_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C81_N30159_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C81_N30159_O_3_C_6_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C89_N30167_O_4_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C89_N30167_O_4_C_5_io_in),
    .io_config(SBMux_C89_N30167_O_4_C_5_io_config),
    .io_out(SBMux_C89_N30167_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C89_N30167_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C89_N30167_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C89_N30167_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C89_N30167_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C97_N30175_O_4_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C97_N30175_O_4_C_5_io_in),
    .io_config(SBMux_C97_N30175_O_4_C_5_io_config),
    .io_out(SBMux_C97_N30175_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C97_N30175_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C97_N30175_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C97_N30175_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C97_N30175_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C1_SCAOptSB SBMux_C101_N30179_O_4_C_1 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C101_N30179_O_4_C_1_io_in),
    .io_config(SBMux_C101_N30179_O_4_C_1_io_config),
    .io_out(SBMux_C101_N30179_O_4_C_1_io_out),
    .io_loopBreak(SBMux_C101_N30179_O_4_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C101_N30179_O_4_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C101_N30179_O_4_C_1_io_cnstClk),
    .io_arst(SBMux_C101_N30179_O_4_C_1_io_arst)
  );
  MuxNInput_O3_C1_SCAOptSB SBMux_C105_N30183_O_3_C_1 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C105_N30183_O_3_C_1_io_in),
    .io_config(SBMux_C105_N30183_O_3_C_1_io_config),
    .io_out(SBMux_C105_N30183_O_3_C_1_io_out),
    .io_loopBreak(SBMux_C105_N30183_O_3_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C105_N30183_O_3_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C105_N30183_O_3_C_1_io_cnstClk),
    .io_arst(SBMux_C105_N30183_O_3_C_1_io_arst)
  );
  MuxNInput_O4_C6_SCAOptSB SBMux_C0_N30186_O_4_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C0_N30186_O_4_C_6_io_in),
    .io_config(SBMux_C0_N30186_O_4_C_6_io_config),
    .io_out(SBMux_C0_N30186_O_4_C_6_io_out),
    .io_loopBreak(SBMux_C0_N30186_O_4_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C0_N30186_O_4_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C0_N30186_O_4_C_6_io_cnstClk),
    .io_arst(SBMux_C0_N30186_O_4_C_6_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C8_N30188_O_4_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C8_N30188_O_4_C_5_io_in),
    .io_config(SBMux_C8_N30188_O_4_C_5_io_config),
    .io_out(SBMux_C8_N30188_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C8_N30188_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C8_N30188_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C8_N30188_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C8_N30188_O_4_C_5_io_arst)
  );
  MuxNInput_O3_C7_SCAOptSB SBMux_C16_N30190_O_3_C_7 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C16_N30190_O_3_C_7_io_in),
    .io_config(SBMux_C16_N30190_O_3_C_7_io_config),
    .io_out(SBMux_C16_N30190_O_3_C_7_io_out),
    .io_loopBreak(SBMux_C16_N30190_O_3_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C16_N30190_O_3_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C16_N30190_O_3_C_7_io_cnstClk),
    .io_arst(SBMux_C16_N30190_O_3_C_7_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C24_N30192_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C24_N30192_O_3_C_6_io_in),
    .io_config(SBMux_C24_N30192_O_3_C_6_io_config),
    .io_out(SBMux_C24_N30192_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C24_N30192_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C24_N30192_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C24_N30192_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C24_N30192_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C32_N30194_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C32_N30194_O_3_C_6_io_in),
    .io_config(SBMux_C32_N30194_O_3_C_6_io_config),
    .io_out(SBMux_C32_N30194_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C32_N30194_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C32_N30194_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C32_N30194_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C32_N30194_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C5_SCAOptSB SBMux_C40_N30196_O_3_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C40_N30196_O_3_C_5_io_in),
    .io_config(SBMux_C40_N30196_O_3_C_5_io_config),
    .io_out(SBMux_C40_N30196_O_3_C_5_io_out),
    .io_loopBreak(SBMux_C40_N30196_O_3_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C40_N30196_O_3_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C40_N30196_O_3_C_5_io_cnstClk),
    .io_arst(SBMux_C40_N30196_O_3_C_5_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C48_N30198_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C48_N30198_O_3_C_6_io_in),
    .io_config(SBMux_C48_N30198_O_3_C_6_io_config),
    .io_out(SBMux_C48_N30198_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C48_N30198_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C48_N30198_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C48_N30198_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C48_N30198_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C56_N30200_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C56_N30200_O_3_C_6_io_in),
    .io_config(SBMux_C56_N30200_O_3_C_6_io_config),
    .io_out(SBMux_C56_N30200_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C56_N30200_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C56_N30200_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C56_N30200_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C56_N30200_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C7_SCAOptSB SBMux_C64_N30202_O_3_C_7 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C64_N30202_O_3_C_7_io_in),
    .io_config(SBMux_C64_N30202_O_3_C_7_io_config),
    .io_out(SBMux_C64_N30202_O_3_C_7_io_out),
    .io_loopBreak(SBMux_C64_N30202_O_3_C_7_io_loopBreak),
    .io_ioGndBle(SBMux_C64_N30202_O_3_C_7_io_ioGndBle),
    .io_cnstClk(SBMux_C64_N30202_O_3_C_7_io_cnstClk),
    .io_arst(SBMux_C64_N30202_O_3_C_7_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C72_N30204_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C72_N30204_O_3_C_6_io_in),
    .io_config(SBMux_C72_N30204_O_3_C_6_io_config),
    .io_out(SBMux_C72_N30204_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C72_N30204_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C72_N30204_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C72_N30204_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C72_N30204_O_3_C_6_io_arst)
  );
  MuxNInput_O3_C6_SCAOptSB SBMux_C80_N30206_O_3_C_6 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C80_N30206_O_3_C_6_io_in),
    .io_config(SBMux_C80_N30206_O_3_C_6_io_config),
    .io_out(SBMux_C80_N30206_O_3_C_6_io_out),
    .io_loopBreak(SBMux_C80_N30206_O_3_C_6_io_loopBreak),
    .io_ioGndBle(SBMux_C80_N30206_O_3_C_6_io_ioGndBle),
    .io_cnstClk(SBMux_C80_N30206_O_3_C_6_io_cnstClk),
    .io_arst(SBMux_C80_N30206_O_3_C_6_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C88_N30208_O_4_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C88_N30208_O_4_C_5_io_in),
    .io_config(SBMux_C88_N30208_O_4_C_5_io_config),
    .io_out(SBMux_C88_N30208_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C88_N30208_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C88_N30208_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C88_N30208_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C88_N30208_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C5_SCAOptSB SBMux_C96_N30210_O_4_C_5 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C96_N30210_O_4_C_5_io_in),
    .io_config(SBMux_C96_N30210_O_4_C_5_io_config),
    .io_out(SBMux_C96_N30210_O_4_C_5_io_out),
    .io_loopBreak(SBMux_C96_N30210_O_4_C_5_io_loopBreak),
    .io_ioGndBle(SBMux_C96_N30210_O_4_C_5_io_ioGndBle),
    .io_cnstClk(SBMux_C96_N30210_O_4_C_5_io_cnstClk),
    .io_arst(SBMux_C96_N30210_O_4_C_5_io_arst)
  );
  MuxNInput_O4_C1_SCAOptSB SBMux_C100_N30212_O_4_C_1 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C100_N30212_O_4_C_1_io_in),
    .io_config(SBMux_C100_N30212_O_4_C_1_io_config),
    .io_out(SBMux_C100_N30212_O_4_C_1_io_out),
    .io_loopBreak(SBMux_C100_N30212_O_4_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C100_N30212_O_4_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C100_N30212_O_4_C_1_io_cnstClk),
    .io_arst(SBMux_C100_N30212_O_4_C_1_io_arst)
  );
  MuxNInput_O3_C1_SCAOptSB SBMux_C104_N30214_O_3_C_1 ( // @[TileFull.scala 141:27]
    .io_in(SBMux_C104_N30214_O_3_C_1_io_in),
    .io_config(SBMux_C104_N30214_O_3_C_1_io_config),
    .io_out(SBMux_C104_N30214_O_3_C_1_io_out),
    .io_loopBreak(SBMux_C104_N30214_O_3_C_1_io_loopBreak),
    .io_ioGndBle(SBMux_C104_N30214_O_3_C_1_io_ioGndBle),
    .io_cnstClk(SBMux_C104_N30214_O_3_C_1_io_cnstClk),
    .io_arst(SBMux_C104_N30214_O_3_C_1_io_arst)
  );
  assign OUT_CHANX_N23695_49 = SBMux_C49_N23695_O_3_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14842_80 = logicBlock_OPIN_80; // @[TileFull.scala 219:12]
  assign OUT_CHANX_N23824_100 = SBMux_C100_N23824_O_0_C_1_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14846_84 = logicBlock_OPIN_84; // @[TileFull.scala 219:12]
  assign OUT_OPIN_N14850_88 = logicBlock_OPIN_88; // @[TileFull.scala 219:12]
  assign OUT_CHANY_N30196_40 = SBMux_C40_N30196_O_3_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23802_16 = SBMux_C16_N23802_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23691_33 = SBMux_C33_N23691_O_3_C_7_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14847_85 = logicBlock_OPIN_85; // @[TileFull.scala 219:12]
  assign OUT_CHANY_N30175_97 = SBMux_C97_N30175_O_4_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30212_100 = SBMux_C100_N30212_O_4_C_1_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23798_0 = SBMux_C0_N23798_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30198_48 = SBMux_C48_N30198_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14840_78 = logicBlock_OPIN_78; // @[TileFull.scala 219:12]
  assign OUT_CHANX_N23685_9 = SBMux_C9_N23685_O_3_C_7_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14844_82 = logicBlock_OPIN_82; // @[TileFull.scala 219:12]
  assign OUT_CHANX_N23816_72 = SBMux_C72_N23816_O_3_C_7_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23769_105 = SBMux_C105_N23769_O_0_C_1_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23683_1 = SBMux_C1_N23683_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23826_104 = SBMux_C104_N23826_O_0_C_1_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23810_48 = SBMux_C48_N23810_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14837_75 = logicBlock_OPIN_75; // @[TileFull.scala 219:12]
  assign OUT_CHANX_N23822_96 = SBMux_C96_N23822_O_2_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30204_72 = SBMux_C72_N30204_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14836_74 = logicBlock_OPIN_74; // @[TileFull.scala 219:12]
  assign OUT_CHANX_N23800_8 = SBMux_C8_N23800_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23804_24 = SBMux_C24_N23804_O_3_C_7_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23812_56 = SBMux_C56_N23812_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14845_83 = logicBlock_OPIN_83; // @[TileFull.scala 219:12]
  assign OUT_CHANY_N30190_16 = SBMux_C16_N30190_O_3_C_7_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30159_81 = SBMux_C81_N30159_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30214_104 = SBMux_C104_N30214_O_3_C_1_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23707_97 = SBMux_C97_N23707_O_2_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14843_81 = logicBlock_OPIN_81; // @[TileFull.scala 219:12]
  assign OUT_CHANX_N23808_40 = SBMux_C40_N23808_O_3_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30087_9 = SBMux_C9_N30087_O_4_C_7_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30206_80 = SBMux_C80_N30206_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30208_88 = SBMux_C88_N30208_O_4_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30119_41 = SBMux_C41_N30119_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14849_87 = logicBlock_OPIN_87; // @[TileFull.scala 219:12]
  assign OUT_CHANY_N30192_24 = SBMux_C24_N30192_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30143_65 = SBMux_C65_N30143_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30095_17 = SBMux_C17_N30095_O_3_C_7_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30186_0 = SBMux_C0_N30186_O_4_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14835_73 = logicBlock_OPIN_73; // @[TileFull.scala 219:12]
  assign OUT_CHANX_N23701_73 = SBMux_C73_N23701_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23689_25 = SBMux_C25_N23689_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23814_64 = SBMux_C64_N23814_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23697_57 = SBMux_C57_N23697_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23687_17 = SBMux_C17_N23687_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30202_64 = SBMux_C64_N30202_O_3_C_7_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14841_79 = logicBlock_OPIN_79; // @[TileFull.scala 219:12]
  assign OUT_OPIN_N14838_76 = logicBlock_OPIN_76; // @[TileFull.scala 219:12]
  assign OUT_CHANX_N23699_65 = SBMux_C65_N23699_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23767_101 = SBMux_C101_N23767_O_0_C_1_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30194_32 = SBMux_C32_N30194_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30188_8 = SBMux_C8_N30188_O_4_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23818_80 = SBMux_C80_N23818_O_2_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30210_96 = SBMux_C96_N30210_O_4_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14839_77 = logicBlock_OPIN_77; // @[TileFull.scala 219:12]
  assign OUT_CHANX_N23703_81 = SBMux_C81_N23703_O_2_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30200_56 = SBMux_C56_N30200_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30167_89 = SBMux_C89_N30167_O_4_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_OPIN_N14848_86 = logicBlock_OPIN_86; // @[TileFull.scala 219:12]
  assign OUT_CHANX_N23693_41 = SBMux_C41_N23693_O_3_C_6_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23820_88 = SBMux_C88_N23820_O_3_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23806_32 = SBMux_C32_N23806_O_3_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30183_105 = SBMux_C105_N30183_O_3_C_1_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANX_N23705_89 = SBMux_C89_N23705_O_3_C_5_io_out; // @[TileFull.scala 146:25]
  assign OUT_CHANY_N30179_101 = SBMux_C101_N30179_O_4_C_1_io_out; // @[TileFull.scala 146:25]
  assign ioConf_confOut = configBlock_ioBundle_confOut[652:0]; // @[TileFull.scala 77:12]
  assign ioConf_scan_out = configBlock_ioBundle_scan_out; // @[TileFull.scala 77:12]
  assign logicBlock_IPIN_0 = CBMux_IPIN0_N14762_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_1 = CBMux_IPIN1_N14763_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_2 = CBMux_IPIN2_N14764_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_3 = CBMux_IPIN3_N14765_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_4 = CBMux_IPIN4_N14766_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_5 = CBMux_IPIN5_N14767_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_6 = CBMux_IPIN6_N14768_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_7 = CBMux_IPIN7_N14769_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_8 = CBMux_IPIN8_N14770_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_9 = CBMux_IPIN9_N14771_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_10 = CBMux_IPIN10_N14772_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_11 = CBMux_IPIN11_N14773_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_12 = CBMux_IPIN12_N14774_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_13 = CBMux_IPIN13_N14775_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_14 = CBMux_IPIN14_N14776_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_15 = CBMux_IPIN15_N14777_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_16 = CBMux_IPIN16_N14778_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_17 = CBMux_IPIN17_N14779_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_18 = CBMux_IPIN18_N14780_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_19 = CBMux_IPIN19_N14781_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_20 = CBMux_IPIN20_N14782_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_21 = CBMux_IPIN21_N14783_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_22 = CBMux_IPIN22_N14784_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_23 = CBMux_IPIN23_N14785_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_24 = CBMux_IPIN24_N14786_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_25 = CBMux_IPIN25_N14787_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_26 = CBMux_IPIN26_N14788_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_27 = CBMux_IPIN27_N14789_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_28 = CBMux_IPIN28_N14790_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_29 = CBMux_IPIN29_N14791_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_30 = CBMux_IPIN30_N14792_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_31 = CBMux_IPIN31_N14793_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_32 = CBMux_IPIN32_N14794_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_33 = CBMux_IPIN33_N14795_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_34 = CBMux_IPIN34_N14796_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_35 = CBMux_IPIN35_N14797_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_36 = CBMux_IPIN36_N14798_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_37 = CBMux_IPIN37_N14799_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_38 = CBMux_IPIN38_N14800_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_39 = CBMux_IPIN39_N14801_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_40 = CBMux_IPIN40_N14802_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_41 = CBMux_IPIN41_N14803_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_42 = CBMux_IPIN42_N14804_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_43 = CBMux_IPIN43_N14805_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_44 = CBMux_IPIN44_N14806_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_45 = CBMux_IPIN45_N14807_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_46 = CBMux_IPIN46_N14808_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_47 = CBMux_IPIN47_N14809_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_48 = CBMux_IPIN48_N14810_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_49 = CBMux_IPIN49_N14811_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_50 = CBMux_IPIN50_N14812_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_51 = CBMux_IPIN51_N14813_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_52 = CBMux_IPIN52_N14814_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_53 = CBMux_IPIN53_N14815_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_54 = CBMux_IPIN54_N14816_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_55 = CBMux_IPIN55_N14817_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_56 = CBMux_IPIN56_N14818_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_57 = CBMux_IPIN57_N14819_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_58 = CBMux_IPIN58_N14820_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_59 = CBMux_IPIN59_N14821_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_60 = CBMux_IPIN60_N14822_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_61 = CBMux_IPIN61_N14823_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_62 = CBMux_IPIN62_N14824_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_63 = CBMux_IPIN63_N14825_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_64 = CBMux_IPIN64_N14826_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_65 = CBMux_IPIN65_N14827_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_66 = CBMux_IPIN66_N14828_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_67 = CBMux_IPIN67_N14829_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_68 = CBMux_IPIN68_N14830_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_69 = CBMux_IPIN69_N14831_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_70 = CBMux_IPIN70_N14832_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_IPIN_71 = CBMux_IPIN71_N14833_io_out; // @[TileFull.scala 106:44]
  assign logicBlock_clock = clock; // @[TileFull.scala 215:26]
  assign logicBlock_reset = reset; // @[TileFull.scala 216:26]
  assign logicBlock_configBits = configBlock_ioBundle_confOut[193:0]; // @[TileFull.scala 214:31]
  assign logicBlock_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 213:30]
  assign logicBlock_gndLBouts = ctrlSignals_gndBlkOuts; // @[TileFull.scala 212:30]
  assign configBlock_clock = ctrlSignals_confClock; // @[TileFull.scala 78:27]
  assign configBlock_ioBundle_scan_in = ioConf_scan_in; // @[TileFull.scala 77:12]
  assign configBlock_ioBundle_scan_en = ioConf_scan_en; // @[TileFull.scala 77:12]
  assign CBMux_IPIN0_N14762_io_in = {CBMux_IPIN0_N14762_io_in_hi,CBMux_IPIN0_N14762_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN0_N14762_io_config = configBlock_ioBundle_confOut[198:194]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN0_N14762_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN0_N14762_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN0_N14762_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN1_N14763_io_in = {CBMux_IPIN1_N14763_io_in_hi,CBMux_IPIN1_N14763_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN1_N14763_io_config = configBlock_ioBundle_confOut[203:199]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN1_N14763_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN1_N14763_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN1_N14763_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN2_N14764_io_in = {CBMux_IPIN2_N14764_io_in_hi,CBMux_IPIN2_N14764_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN2_N14764_io_config = configBlock_ioBundle_confOut[208:204]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN2_N14764_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN2_N14764_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN2_N14764_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN3_N14765_io_in = {CBMux_IPIN3_N14765_io_in_hi,CBMux_IPIN3_N14765_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN3_N14765_io_config = configBlock_ioBundle_confOut[213:209]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN3_N14765_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN3_N14765_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN3_N14765_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN4_N14766_io_in = {CBMux_IPIN4_N14766_io_in_hi,CBMux_IPIN4_N14766_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN4_N14766_io_config = configBlock_ioBundle_confOut[218:214]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN4_N14766_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN4_N14766_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN4_N14766_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN5_N14767_io_in = {CBMux_IPIN5_N14767_io_in_hi,CBMux_IPIN5_N14767_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN5_N14767_io_config = configBlock_ioBundle_confOut[223:219]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN5_N14767_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN5_N14767_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN5_N14767_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN6_N14768_io_in = {CBMux_IPIN6_N14768_io_in_hi,CBMux_IPIN6_N14768_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN6_N14768_io_config = configBlock_ioBundle_confOut[228:224]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN6_N14768_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN6_N14768_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN6_N14768_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN7_N14769_io_in = {CBMux_IPIN7_N14769_io_in_hi,CBMux_IPIN7_N14769_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN7_N14769_io_config = configBlock_ioBundle_confOut[233:229]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN7_N14769_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN7_N14769_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN7_N14769_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN8_N14770_io_in = {CBMux_IPIN7_N14769_io_in_hi,CBMux_IPIN8_N14770_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN8_N14770_io_config = configBlock_ioBundle_confOut[238:234]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN8_N14770_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN8_N14770_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN8_N14770_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN9_N14771_io_in = {CBMux_IPIN9_N14771_io_in_hi,CBMux_IPIN9_N14771_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN9_N14771_io_config = configBlock_ioBundle_confOut[243:239]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN9_N14771_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN9_N14771_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN9_N14771_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN10_N14772_io_in = {CBMux_IPIN10_N14772_io_in_hi,CBMux_IPIN10_N14772_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN10_N14772_io_config = configBlock_ioBundle_confOut[248:244]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN10_N14772_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN10_N14772_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN10_N14772_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN11_N14773_io_in = {CBMux_IPIN6_N14768_io_in_hi,CBMux_IPIN11_N14773_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN11_N14773_io_config = configBlock_ioBundle_confOut[253:249]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN11_N14773_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN11_N14773_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN11_N14773_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN12_N14774_io_in = {CBMux_IPIN12_N14774_io_in_hi,CBMux_IPIN12_N14774_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN12_N14774_io_config = configBlock_ioBundle_confOut[258:254]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN12_N14774_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN12_N14774_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN12_N14774_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN13_N14775_io_in = {CBMux_IPIN13_N14775_io_in_hi,CBMux_IPIN13_N14775_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN13_N14775_io_config = configBlock_ioBundle_confOut[263:259]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN13_N14775_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN13_N14775_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN13_N14775_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN14_N14776_io_in = {CBMux_IPIN14_N14776_io_in_hi,CBMux_IPIN14_N14776_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN14_N14776_io_config = configBlock_ioBundle_confOut[268:264]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN14_N14776_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN14_N14776_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN14_N14776_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN15_N14777_io_in = {CBMux_IPIN15_N14777_io_in_hi,CBMux_IPIN15_N14777_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN15_N14777_io_config = configBlock_ioBundle_confOut[273:269]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN15_N14777_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN15_N14777_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN15_N14777_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN16_N14778_io_in = {CBMux_IPIN16_N14778_io_in_hi,CBMux_IPIN16_N14778_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN16_N14778_io_config = configBlock_ioBundle_confOut[278:274]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN16_N14778_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN16_N14778_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN16_N14778_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN17_N14779_io_in = {CBMux_IPIN17_N14779_io_in_hi,CBMux_IPIN17_N14779_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN17_N14779_io_config = configBlock_ioBundle_confOut[283:279]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN17_N14779_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN17_N14779_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN17_N14779_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN18_N14780_io_in = {CBMux_IPIN18_N14780_io_in_hi,CBMux_IPIN18_N14780_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN18_N14780_io_config = configBlock_ioBundle_confOut[288:284]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN18_N14780_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN18_N14780_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN18_N14780_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN19_N14781_io_in = {CBMux_IPIN19_N14781_io_in_hi,CBMux_IPIN19_N14781_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN19_N14781_io_config = configBlock_ioBundle_confOut[293:289]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN19_N14781_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN19_N14781_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN19_N14781_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN20_N14782_io_in = {CBMux_IPIN20_N14782_io_in_hi,CBMux_IPIN20_N14782_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN20_N14782_io_config = configBlock_ioBundle_confOut[298:294]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN20_N14782_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN20_N14782_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN20_N14782_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN21_N14783_io_in = {CBMux_IPIN21_N14783_io_in_hi,CBMux_IPIN21_N14783_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN21_N14783_io_config = configBlock_ioBundle_confOut[303:299]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN21_N14783_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN21_N14783_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN21_N14783_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN22_N14784_io_in = {CBMux_IPIN22_N14784_io_in_hi,CBMux_IPIN22_N14784_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN22_N14784_io_config = configBlock_ioBundle_confOut[308:304]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN22_N14784_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN22_N14784_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN22_N14784_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN23_N14785_io_in = {CBMux_IPIN23_N14785_io_in_hi,CBMux_IPIN23_N14785_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN23_N14785_io_config = configBlock_ioBundle_confOut[313:309]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN23_N14785_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN23_N14785_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN23_N14785_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN24_N14786_io_in = {CBMux_IPIN24_N14786_io_in_hi,CBMux_IPIN24_N14786_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN24_N14786_io_config = configBlock_ioBundle_confOut[318:314]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN24_N14786_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN24_N14786_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN24_N14786_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN25_N14787_io_in = {CBMux_IPIN25_N14787_io_in_hi,CBMux_IPIN25_N14787_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN25_N14787_io_config = configBlock_ioBundle_confOut[323:319]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN25_N14787_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN25_N14787_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN25_N14787_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN26_N14788_io_in = {CBMux_IPIN26_N14788_io_in_hi,CBMux_IPIN26_N14788_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN26_N14788_io_config = configBlock_ioBundle_confOut[328:324]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN26_N14788_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN26_N14788_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN26_N14788_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN27_N14789_io_in = {CBMux_IPIN27_N14789_io_in_hi,CBMux_IPIN27_N14789_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN27_N14789_io_config = configBlock_ioBundle_confOut[333:329]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN27_N14789_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN27_N14789_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN27_N14789_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN28_N14790_io_in = {CBMux_IPIN28_N14790_io_in_hi,CBMux_IPIN28_N14790_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN28_N14790_io_config = configBlock_ioBundle_confOut[338:334]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN28_N14790_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN28_N14790_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN28_N14790_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN29_N14791_io_in = {CBMux_IPIN29_N14791_io_in_hi,CBMux_IPIN29_N14791_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN29_N14791_io_config = configBlock_ioBundle_confOut[343:339]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN29_N14791_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN29_N14791_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN29_N14791_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN30_N14792_io_in = {CBMux_IPIN30_N14792_io_in_hi,CBMux_IPIN30_N14792_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN30_N14792_io_config = configBlock_ioBundle_confOut[348:344]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN30_N14792_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN30_N14792_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN30_N14792_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN31_N14793_io_in = {CBMux_IPIN26_N14788_io_in_hi,CBMux_IPIN26_N14788_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN31_N14793_io_config = configBlock_ioBundle_confOut[353:349]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN31_N14793_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN31_N14793_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN31_N14793_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN32_N14794_io_in = {CBMux_IPIN32_N14794_io_in_hi,CBMux_IPIN32_N14794_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN32_N14794_io_config = configBlock_ioBundle_confOut[358:354]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN32_N14794_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN32_N14794_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN32_N14794_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN33_N14795_io_in = {CBMux_IPIN33_N14795_io_in_hi,CBMux_IPIN33_N14795_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN33_N14795_io_config = configBlock_ioBundle_confOut[363:359]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN33_N14795_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN33_N14795_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN33_N14795_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN34_N14796_io_in = {CBMux_IPIN25_N14787_io_in_hi,CBMux_IPIN25_N14787_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN34_N14796_io_config = configBlock_ioBundle_confOut[368:364]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN34_N14796_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN34_N14796_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN34_N14796_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN35_N14797_io_in = {CBMux_IPIN35_N14797_io_in_hi,CBMux_IPIN35_N14797_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN35_N14797_io_config = configBlock_ioBundle_confOut[373:369]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN35_N14797_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN35_N14797_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN35_N14797_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN36_N14798_io_in = {CBMux_IPIN36_N14798_io_in_hi,CBMux_IPIN36_N14798_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN36_N14798_io_config = configBlock_ioBundle_confOut[378:374]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN36_N14798_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN36_N14798_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN36_N14798_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN37_N14799_io_in = {CBMux_IPIN37_N14799_io_in_hi,CBMux_IPIN37_N14799_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN37_N14799_io_config = configBlock_ioBundle_confOut[383:379]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN37_N14799_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN37_N14799_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN37_N14799_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN38_N14800_io_in = {CBMux_IPIN38_N14800_io_in_hi,CBMux_IPIN38_N14800_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN38_N14800_io_config = configBlock_ioBundle_confOut[388:384]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN38_N14800_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN38_N14800_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN38_N14800_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN39_N14801_io_in = {CBMux_IPIN39_N14801_io_in_hi,CBMux_IPIN39_N14801_io_in_lo}; // @[TileFull.scala 175:8]
  assign CBMux_IPIN39_N14801_io_config = configBlock_ioBundle_confOut[393:389]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN39_N14801_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN39_N14801_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN39_N14801_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN40_N14802_io_in = IN_OPIN_N15095_89; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN40_N14802_io_config = configBlock_ioBundle_confOut[394]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN40_N14802_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN40_N14802_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN40_N14802_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN41_N14803_io_in = IN_OPIN_N15096_90; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN41_N14803_io_config = configBlock_ioBundle_confOut[395]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN41_N14803_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN41_N14803_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN41_N14803_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN42_N14804_io_in = IN_OPIN_N15097_91; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN42_N14804_io_config = configBlock_ioBundle_confOut[396]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN42_N14804_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN42_N14804_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN42_N14804_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN43_N14805_io_in = IN_OPIN_N15098_92; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN43_N14805_io_config = configBlock_ioBundle_confOut[397]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN43_N14805_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN43_N14805_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN43_N14805_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN44_N14806_io_in = IN_OPIN_N15099_93; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN44_N14806_io_config = configBlock_ioBundle_confOut[398]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN44_N14806_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN44_N14806_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN44_N14806_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN45_N14807_io_in = IN_OPIN_N15100_94; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN45_N14807_io_config = configBlock_ioBundle_confOut[399]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN45_N14807_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN45_N14807_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN45_N14807_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN46_N14808_io_in = IN_OPIN_N15101_95; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN46_N14808_io_config = configBlock_ioBundle_confOut[400]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN46_N14808_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN46_N14808_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN46_N14808_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN47_N14809_io_in = IN_OPIN_N15102_96; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN47_N14809_io_config = configBlock_ioBundle_confOut[401]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN47_N14809_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN47_N14809_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN47_N14809_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN48_N14810_io_in = IN_OPIN_N15103_97; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN48_N14810_io_config = configBlock_ioBundle_confOut[402]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN48_N14810_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN48_N14810_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN48_N14810_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN49_N14811_io_in = IN_OPIN_N15104_98; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN49_N14811_io_config = configBlock_ioBundle_confOut[403]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN49_N14811_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN49_N14811_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN49_N14811_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN50_N14812_io_in = IN_OPIN_N15105_99; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN50_N14812_io_config = configBlock_ioBundle_confOut[404]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN50_N14812_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN50_N14812_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN50_N14812_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN51_N14813_io_in = IN_OPIN_N15106_100; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN51_N14813_io_config = configBlock_ioBundle_confOut[405]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN51_N14813_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN51_N14813_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN51_N14813_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN52_N14814_io_in = IN_OPIN_N15107_101; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN52_N14814_io_config = configBlock_ioBundle_confOut[406]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN52_N14814_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN52_N14814_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN52_N14814_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN53_N14815_io_in = IN_OPIN_N15108_102; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN53_N14815_io_config = configBlock_ioBundle_confOut[407]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN53_N14815_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN53_N14815_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN53_N14815_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN54_N14816_io_in = IN_OPIN_N15109_103; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN54_N14816_io_config = configBlock_ioBundle_confOut[408]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN54_N14816_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN54_N14816_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN54_N14816_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN55_N14817_io_in = IN_OPIN_N15110_104; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN55_N14817_io_config = configBlock_ioBundle_confOut[409]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN55_N14817_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN55_N14817_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN55_N14817_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN56_N14818_io_in = IN_OPIN_N15111_105; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN56_N14818_io_config = configBlock_ioBundle_confOut[410]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN56_N14818_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN56_N14818_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN56_N14818_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN57_N14819_io_in = IN_OPIN_N15112_106; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN57_N14819_io_config = configBlock_ioBundle_confOut[411]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN57_N14819_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN57_N14819_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN57_N14819_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN58_N14820_io_in = IN_OPIN_N15113_107; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN58_N14820_io_config = configBlock_ioBundle_confOut[412]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN58_N14820_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN58_N14820_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN58_N14820_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN59_N14821_io_in = IN_OPIN_N15114_108; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN59_N14821_io_config = configBlock_ioBundle_confOut[413]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN59_N14821_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN59_N14821_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN59_N14821_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN60_N14822_io_in = IN_OPIN_N15115_109; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN60_N14822_io_config = configBlock_ioBundle_confOut[414]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN60_N14822_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN60_N14822_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN60_N14822_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN61_N14823_io_in = IN_OPIN_N15116_110; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN61_N14823_io_config = configBlock_ioBundle_confOut[415]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN61_N14823_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN61_N14823_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN61_N14823_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN62_N14824_io_in = IN_OPIN_N15117_111; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN62_N14824_io_config = configBlock_ioBundle_confOut[416]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN62_N14824_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN62_N14824_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN62_N14824_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN63_N14825_io_in = IN_OPIN_N15118_112; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN63_N14825_io_config = configBlock_ioBundle_confOut[417]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN63_N14825_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN63_N14825_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN63_N14825_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN64_N14826_io_in = IN_OPIN_N15119_113; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN64_N14826_io_config = configBlock_ioBundle_confOut[418]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN64_N14826_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN64_N14826_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN64_N14826_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN65_N14827_io_in = IN_OPIN_N15120_114; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN65_N14827_io_config = configBlock_ioBundle_confOut[419]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN65_N14827_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN65_N14827_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN65_N14827_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN66_N14828_io_in = IN_OPIN_N15121_115; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN66_N14828_io_config = configBlock_ioBundle_confOut[420]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN66_N14828_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN66_N14828_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN66_N14828_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN67_N14829_io_in = IN_OPIN_N15122_116; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN67_N14829_io_config = configBlock_ioBundle_confOut[421]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN67_N14829_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN67_N14829_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN67_N14829_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN68_N14830_io_in = IN_OPIN_N15123_117; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN68_N14830_io_config = configBlock_ioBundle_confOut[422]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN68_N14830_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN68_N14830_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN68_N14830_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN69_N14831_io_in = IN_OPIN_N15124_118; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN69_N14831_io_config = configBlock_ioBundle_confOut[423]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN69_N14831_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN69_N14831_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN69_N14831_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN70_N14832_io_in = IN_OPIN_N15125_119; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN70_N14832_io_config = configBlock_ioBundle_confOut[424]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN70_N14832_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN70_N14832_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN70_N14832_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign CBMux_IPIN71_N14833_io_in = IN_OPIN_N15126_120; // @[TileFull.scala 170:{37,37}]
  assign CBMux_IPIN71_N14833_io_config = configBlock_ioBundle_confOut[425]; // @[TileFull.scala 110:62]
  assign CBMux_IPIN71_N14833_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 113:30]
  assign CBMux_IPIN71_N14833_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 114:28]
  assign CBMux_IPIN71_N14833_io_arst = ctrlSignals_arst; // @[TileFull.scala 115:25]
  assign SBMux_C1_N23683_O_3_C_6_io_in = {SBMux_C1_N23683_O_3_C_6_io_in_hi,SBMux_C1_N23683_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C1_N23683_O_3_C_6_io_config = configBlock_ioBundle_confOut[429:426]; // @[TileFull.scala 151:60]
  assign SBMux_C1_N23683_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C1_N23683_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C1_N23683_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C1_N23683_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C9_N23685_O_3_C_7_io_in = {SBMux_C9_N23685_O_3_C_7_io_in_hi,SBMux_C9_N23685_O_3_C_7_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C9_N23685_O_3_C_7_io_config = configBlock_ioBundle_confOut[433:430]; // @[TileFull.scala 151:60]
  assign SBMux_C9_N23685_O_3_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C9_N23685_O_3_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C9_N23685_O_3_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C9_N23685_O_3_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C17_N23687_O_3_C_6_io_in = {SBMux_C17_N23687_O_3_C_6_io_in_hi,SBMux_C17_N23687_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C17_N23687_O_3_C_6_io_config = configBlock_ioBundle_confOut[437:434]; // @[TileFull.scala 151:60]
  assign SBMux_C17_N23687_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C17_N23687_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C17_N23687_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C17_N23687_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C25_N23689_O_3_C_6_io_in = {SBMux_C25_N23689_O_3_C_6_io_in_hi,SBMux_C25_N23689_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C25_N23689_O_3_C_6_io_config = configBlock_ioBundle_confOut[441:438]; // @[TileFull.scala 151:60]
  assign SBMux_C25_N23689_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C25_N23689_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C25_N23689_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C25_N23689_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C33_N23691_O_3_C_7_io_in = {SBMux_C33_N23691_O_3_C_7_io_in_hi,SBMux_C33_N23691_O_3_C_7_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C33_N23691_O_3_C_7_io_config = configBlock_ioBundle_confOut[445:442]; // @[TileFull.scala 151:60]
  assign SBMux_C33_N23691_O_3_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C33_N23691_O_3_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C33_N23691_O_3_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C33_N23691_O_3_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C41_N23693_O_3_C_6_io_in = {SBMux_C41_N23693_O_3_C_6_io_in_hi,SBMux_C41_N23693_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C41_N23693_O_3_C_6_io_config = configBlock_ioBundle_confOut[449:446]; // @[TileFull.scala 151:60]
  assign SBMux_C41_N23693_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C41_N23693_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C41_N23693_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C41_N23693_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C49_N23695_O_3_C_5_io_in = {SBMux_C49_N23695_O_3_C_5_io_in_hi,SBMux_C49_N23695_O_3_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C49_N23695_O_3_C_5_io_config = configBlock_ioBundle_confOut[453:450]; // @[TileFull.scala 151:60]
  assign SBMux_C49_N23695_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C49_N23695_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C49_N23695_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C49_N23695_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C57_N23697_O_3_C_6_io_in = {SBMux_C57_N23697_O_3_C_6_io_in_hi,SBMux_C57_N23697_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C57_N23697_O_3_C_6_io_config = configBlock_ioBundle_confOut[457:454]; // @[TileFull.scala 151:60]
  assign SBMux_C57_N23697_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C57_N23697_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C57_N23697_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C57_N23697_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C65_N23699_O_3_C_6_io_in = {SBMux_C65_N23699_O_3_C_6_io_in_hi,SBMux_C65_N23699_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C65_N23699_O_3_C_6_io_config = configBlock_ioBundle_confOut[461:458]; // @[TileFull.scala 151:60]
  assign SBMux_C65_N23699_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C65_N23699_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C65_N23699_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C65_N23699_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C73_N23701_O_3_C_6_io_in = {SBMux_C73_N23701_O_3_C_6_io_in_hi,SBMux_C73_N23701_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C73_N23701_O_3_C_6_io_config = configBlock_ioBundle_confOut[465:462]; // @[TileFull.scala 151:60]
  assign SBMux_C73_N23701_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C73_N23701_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C73_N23701_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C73_N23701_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C81_N23703_O_2_C_5_io_in = {SBMux_C81_N23703_O_2_C_5_io_in_hi,SBMux_C81_N23703_O_2_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C81_N23703_O_2_C_5_io_config = configBlock_ioBundle_confOut[469:466]; // @[TileFull.scala 151:60]
  assign SBMux_C81_N23703_O_2_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C81_N23703_O_2_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C81_N23703_O_2_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C81_N23703_O_2_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C89_N23705_O_3_C_5_io_in = {SBMux_C89_N23705_O_3_C_5_io_in_hi,SBMux_C89_N23705_O_3_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C89_N23705_O_3_C_5_io_config = configBlock_ioBundle_confOut[473:470]; // @[TileFull.scala 151:60]
  assign SBMux_C89_N23705_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C89_N23705_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C89_N23705_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C89_N23705_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C97_N23707_O_2_C_5_io_in = {SBMux_C97_N23707_O_2_C_5_io_in_hi,SBMux_C97_N23707_O_2_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C97_N23707_O_2_C_5_io_config = configBlock_ioBundle_confOut[477:474]; // @[TileFull.scala 151:60]
  assign SBMux_C97_N23707_O_2_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C97_N23707_O_2_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C97_N23707_O_2_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C97_N23707_O_2_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C101_N23767_O_0_C_1_io_in = IN_CHANX_N23827_105; // @[TileFull.scala 187:{39,39}]
  assign SBMux_C101_N23767_O_0_C_1_io_config = configBlock_ioBundle_confOut[479:478]; // @[TileFull.scala 151:60]
  assign SBMux_C101_N23767_O_0_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C101_N23767_O_0_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C101_N23767_O_0_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C101_N23767_O_0_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C105_N23769_O_0_C_1_io_in = IN_CHANX_N23825_101; // @[TileFull.scala 187:{39,39}]
  assign SBMux_C105_N23769_O_0_C_1_io_config = configBlock_ioBundle_confOut[481:480]; // @[TileFull.scala 151:60]
  assign SBMux_C105_N23769_O_0_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C105_N23769_O_0_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C105_N23769_O_0_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C105_N23769_O_0_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C0_N23798_O_3_C_6_io_in = {SBMux_C0_N23798_O_3_C_6_io_in_hi,SBMux_C0_N23798_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C0_N23798_O_3_C_6_io_config = configBlock_ioBundle_confOut[485:482]; // @[TileFull.scala 151:60]
  assign SBMux_C0_N23798_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C0_N23798_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C0_N23798_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C0_N23798_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C8_N23800_O_3_C_6_io_in = {SBMux_C8_N23800_O_3_C_6_io_in_hi,SBMux_C8_N23800_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C8_N23800_O_3_C_6_io_config = configBlock_ioBundle_confOut[489:486]; // @[TileFull.scala 151:60]
  assign SBMux_C8_N23800_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C8_N23800_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C8_N23800_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C8_N23800_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C16_N23802_O_3_C_6_io_in = {SBMux_C16_N23802_O_3_C_6_io_in_hi,SBMux_C16_N23802_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C16_N23802_O_3_C_6_io_config = configBlock_ioBundle_confOut[493:490]; // @[TileFull.scala 151:60]
  assign SBMux_C16_N23802_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C16_N23802_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C16_N23802_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C16_N23802_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C24_N23804_O_3_C_7_io_in = {SBMux_C24_N23804_O_3_C_7_io_in_hi,SBMux_C24_N23804_O_3_C_7_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C24_N23804_O_3_C_7_io_config = configBlock_ioBundle_confOut[497:494]; // @[TileFull.scala 151:60]
  assign SBMux_C24_N23804_O_3_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C24_N23804_O_3_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C24_N23804_O_3_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C24_N23804_O_3_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C32_N23806_O_3_C_5_io_in = {SBMux_C32_N23806_O_3_C_5_io_in_hi,SBMux_C32_N23806_O_3_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C32_N23806_O_3_C_5_io_config = configBlock_ioBundle_confOut[501:498]; // @[TileFull.scala 151:60]
  assign SBMux_C32_N23806_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C32_N23806_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C32_N23806_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C32_N23806_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C40_N23808_O_3_C_5_io_in = {SBMux_C40_N23808_O_3_C_5_io_in_hi,SBMux_C40_N23808_O_3_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C40_N23808_O_3_C_5_io_config = configBlock_ioBundle_confOut[505:502]; // @[TileFull.scala 151:60]
  assign SBMux_C40_N23808_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C40_N23808_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C40_N23808_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C40_N23808_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C48_N23810_O_3_C_6_io_in = {SBMux_C48_N23810_O_3_C_6_io_in_hi,SBMux_C48_N23810_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C48_N23810_O_3_C_6_io_config = configBlock_ioBundle_confOut[509:506]; // @[TileFull.scala 151:60]
  assign SBMux_C48_N23810_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C48_N23810_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C48_N23810_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C48_N23810_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C56_N23812_O_3_C_6_io_in = {SBMux_C56_N23812_O_3_C_6_io_in_hi,SBMux_C56_N23812_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C56_N23812_O_3_C_6_io_config = configBlock_ioBundle_confOut[513:510]; // @[TileFull.scala 151:60]
  assign SBMux_C56_N23812_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C56_N23812_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C56_N23812_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C56_N23812_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C64_N23814_O_3_C_6_io_in = {SBMux_C64_N23814_O_3_C_6_io_in_hi,SBMux_C64_N23814_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C64_N23814_O_3_C_6_io_config = configBlock_ioBundle_confOut[517:514]; // @[TileFull.scala 151:60]
  assign SBMux_C64_N23814_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C64_N23814_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C64_N23814_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C64_N23814_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C72_N23816_O_3_C_7_io_in = {SBMux_C72_N23816_O_3_C_7_io_in_hi,SBMux_C72_N23816_O_3_C_7_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C72_N23816_O_3_C_7_io_config = configBlock_ioBundle_confOut[521:518]; // @[TileFull.scala 151:60]
  assign SBMux_C72_N23816_O_3_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C72_N23816_O_3_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C72_N23816_O_3_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C72_N23816_O_3_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C80_N23818_O_2_C_6_io_in = {SBMux_C80_N23818_O_2_C_6_io_in_hi,SBMux_C80_N23818_O_2_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C80_N23818_O_2_C_6_io_config = configBlock_ioBundle_confOut[525:522]; // @[TileFull.scala 151:60]
  assign SBMux_C80_N23818_O_2_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C80_N23818_O_2_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C80_N23818_O_2_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C80_N23818_O_2_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C88_N23820_O_3_C_5_io_in = {SBMux_C88_N23820_O_3_C_5_io_in_hi,SBMux_C88_N23820_O_3_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C88_N23820_O_3_C_5_io_config = configBlock_ioBundle_confOut[529:526]; // @[TileFull.scala 151:60]
  assign SBMux_C88_N23820_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C88_N23820_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C88_N23820_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C88_N23820_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C96_N23822_O_2_C_5_io_in = {SBMux_C96_N23822_O_2_C_5_io_in_hi,SBMux_C96_N23822_O_2_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C96_N23822_O_2_C_5_io_config = configBlock_ioBundle_confOut[533:530]; // @[TileFull.scala 151:60]
  assign SBMux_C96_N23822_O_2_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C96_N23822_O_2_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C96_N23822_O_2_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C96_N23822_O_2_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C100_N23824_O_0_C_1_io_in = IN_CHANX_N23766_100; // @[TileFull.scala 187:{39,39}]
  assign SBMux_C100_N23824_O_0_C_1_io_config = configBlock_ioBundle_confOut[535:534]; // @[TileFull.scala 151:60]
  assign SBMux_C100_N23824_O_0_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C100_N23824_O_0_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C100_N23824_O_0_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C100_N23824_O_0_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C104_N23826_O_0_C_1_io_in = IN_CHANX_N23768_104; // @[TileFull.scala 187:{39,39}]
  assign SBMux_C104_N23826_O_0_C_1_io_config = configBlock_ioBundle_confOut[537:536]; // @[TileFull.scala 151:60]
  assign SBMux_C104_N23826_O_0_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C104_N23826_O_0_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C104_N23826_O_0_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C104_N23826_O_0_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C1_N30079_O_4_C_6_io_in = {SBMux_C1_N30079_O_4_C_6_io_in_hi,SBMux_C1_N30079_O_4_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C1_N30079_O_4_C_6_io_config = configBlock_ioBundle_confOut[541:538]; // @[TileFull.scala 151:60]
  assign SBMux_C1_N30079_O_4_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C1_N30079_O_4_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C1_N30079_O_4_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C1_N30079_O_4_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C9_N30087_O_4_C_7_io_in = {SBMux_C9_N30087_O_4_C_7_io_in_hi,SBMux_C9_N30087_O_4_C_7_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C9_N30087_O_4_C_7_io_config = configBlock_ioBundle_confOut[545:542]; // @[TileFull.scala 151:60]
  assign SBMux_C9_N30087_O_4_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C9_N30087_O_4_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C9_N30087_O_4_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C9_N30087_O_4_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C17_N30095_O_3_C_7_io_in = {SBMux_C17_N30095_O_3_C_7_io_in_hi,SBMux_C17_N30095_O_3_C_7_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C17_N30095_O_3_C_7_io_config = configBlock_ioBundle_confOut[549:546]; // @[TileFull.scala 151:60]
  assign SBMux_C17_N30095_O_3_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C17_N30095_O_3_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C17_N30095_O_3_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C17_N30095_O_3_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C25_N30103_O_3_C_6_io_in = {SBMux_C25_N30103_O_3_C_6_io_in_hi,SBMux_C25_N30103_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C25_N30103_O_3_C_6_io_config = configBlock_ioBundle_confOut[553:550]; // @[TileFull.scala 151:60]
  assign SBMux_C25_N30103_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C25_N30103_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C25_N30103_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C25_N30103_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C33_N30111_O_3_C_4_io_in = {SBMux_C33_N30111_O_3_C_4_io_in_hi,SBMux_C33_N30111_O_3_C_4_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C33_N30111_O_3_C_4_io_config = configBlock_ioBundle_confOut[556:554]; // @[TileFull.scala 151:60]
  assign SBMux_C33_N30111_O_3_C_4_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C33_N30111_O_3_C_4_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C33_N30111_O_3_C_4_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C33_N30111_O_3_C_4_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C41_N30119_O_3_C_6_io_in = {SBMux_C41_N30119_O_3_C_6_io_in_hi,SBMux_C41_N30119_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C41_N30119_O_3_C_6_io_config = configBlock_ioBundle_confOut[560:557]; // @[TileFull.scala 151:60]
  assign SBMux_C41_N30119_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C41_N30119_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C41_N30119_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C41_N30119_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C49_N30127_O_3_C_6_io_in = {SBMux_C49_N30127_O_3_C_6_io_in_hi,SBMux_C41_N30119_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C49_N30127_O_3_C_6_io_config = configBlock_ioBundle_confOut[564:561]; // @[TileFull.scala 151:60]
  assign SBMux_C49_N30127_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C49_N30127_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C49_N30127_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C49_N30127_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C57_N30135_O_3_C_6_io_in = {SBMux_C57_N30135_O_3_C_6_io_in_hi,SBMux_C57_N30135_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C57_N30135_O_3_C_6_io_config = configBlock_ioBundle_confOut[568:565]; // @[TileFull.scala 151:60]
  assign SBMux_C57_N30135_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C57_N30135_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C57_N30135_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C57_N30135_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C65_N30143_O_3_C_6_io_in = {SBMux_C65_N30143_O_3_C_6_io_in_hi,SBMux_C65_N30143_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C65_N30143_O_3_C_6_io_config = configBlock_ioBundle_confOut[572:569]; // @[TileFull.scala 151:60]
  assign SBMux_C65_N30143_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C65_N30143_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C65_N30143_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C65_N30143_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C73_N30151_O_3_C_6_io_in = {SBMux_C73_N30151_O_3_C_6_io_in_hi,SBMux_C73_N30151_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C73_N30151_O_3_C_6_io_config = configBlock_ioBundle_confOut[576:573]; // @[TileFull.scala 151:60]
  assign SBMux_C73_N30151_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C73_N30151_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C73_N30151_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C73_N30151_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C81_N30159_O_3_C_6_io_in = {SBMux_C81_N30159_O_3_C_6_io_in_hi,SBMux_C81_N30159_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C81_N30159_O_3_C_6_io_config = configBlock_ioBundle_confOut[580:577]; // @[TileFull.scala 151:60]
  assign SBMux_C81_N30159_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C81_N30159_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C81_N30159_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C81_N30159_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C89_N30167_O_4_C_5_io_in = {SBMux_C89_N30167_O_4_C_5_io_in_hi,SBMux_C89_N30167_O_4_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C89_N30167_O_4_C_5_io_config = configBlock_ioBundle_confOut[584:581]; // @[TileFull.scala 151:60]
  assign SBMux_C89_N30167_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C89_N30167_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C89_N30167_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C89_N30167_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C97_N30175_O_4_C_5_io_in = {SBMux_C97_N30175_O_4_C_5_io_in_hi,SBMux_C97_N30175_O_4_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C97_N30175_O_4_C_5_io_config = configBlock_ioBundle_confOut[588:585]; // @[TileFull.scala 151:60]
  assign SBMux_C97_N30175_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C97_N30175_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C97_N30175_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C97_N30175_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C101_N30179_O_4_C_1_io_in = {SBMux_C101_N30179_O_4_C_1_io_in_hi,SBMux_C1_N30079_O_4_C_6_io_in_lo_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C101_N30179_O_4_C_1_io_config = configBlock_ioBundle_confOut[591:589]; // @[TileFull.scala 151:60]
  assign SBMux_C101_N30179_O_4_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C101_N30179_O_4_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C101_N30179_O_4_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C101_N30179_O_4_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C105_N30183_O_3_C_1_io_in = {SBMux_C105_N30183_O_3_C_1_io_in_hi,SBMux_C41_N30119_O_3_C_6_io_in_lo_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C105_N30183_O_3_C_1_io_config = configBlock_ioBundle_confOut[594:592]; // @[TileFull.scala 151:60]
  assign SBMux_C105_N30183_O_3_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C105_N30183_O_3_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C105_N30183_O_3_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C105_N30183_O_3_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C0_N30186_O_4_C_6_io_in = {SBMux_C0_N30186_O_4_C_6_io_in_hi,SBMux_C0_N30186_O_4_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C0_N30186_O_4_C_6_io_config = configBlock_ioBundle_confOut[598:595]; // @[TileFull.scala 151:60]
  assign SBMux_C0_N30186_O_4_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C0_N30186_O_4_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C0_N30186_O_4_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C0_N30186_O_4_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C8_N30188_O_4_C_5_io_in = {SBMux_C8_N30188_O_4_C_5_io_in_hi,SBMux_C8_N30188_O_4_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C8_N30188_O_4_C_5_io_config = configBlock_ioBundle_confOut[602:599]; // @[TileFull.scala 151:60]
  assign SBMux_C8_N30188_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C8_N30188_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C8_N30188_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C8_N30188_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C16_N30190_O_3_C_7_io_in = {SBMux_C16_N30190_O_3_C_7_io_in_hi,SBMux_C16_N30190_O_3_C_7_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C16_N30190_O_3_C_7_io_config = configBlock_ioBundle_confOut[606:603]; // @[TileFull.scala 151:60]
  assign SBMux_C16_N30190_O_3_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C16_N30190_O_3_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C16_N30190_O_3_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C16_N30190_O_3_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C24_N30192_O_3_C_6_io_in = {SBMux_C24_N30192_O_3_C_6_io_in_hi,SBMux_C24_N30192_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C24_N30192_O_3_C_6_io_config = configBlock_ioBundle_confOut[610:607]; // @[TileFull.scala 151:60]
  assign SBMux_C24_N30192_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C24_N30192_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C24_N30192_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C24_N30192_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C32_N30194_O_3_C_6_io_in = {SBMux_C32_N30194_O_3_C_6_io_in_hi,SBMux_C32_N30194_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C32_N30194_O_3_C_6_io_config = configBlock_ioBundle_confOut[614:611]; // @[TileFull.scala 151:60]
  assign SBMux_C32_N30194_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C32_N30194_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C32_N30194_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C32_N30194_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C40_N30196_O_3_C_5_io_in = {SBMux_C40_N30196_O_3_C_5_io_in_hi,SBMux_C40_N30196_O_3_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C40_N30196_O_3_C_5_io_config = configBlock_ioBundle_confOut[618:615]; // @[TileFull.scala 151:60]
  assign SBMux_C40_N30196_O_3_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C40_N30196_O_3_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C40_N30196_O_3_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C40_N30196_O_3_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C48_N30198_O_3_C_6_io_in = {SBMux_C48_N30198_O_3_C_6_io_in_hi,SBMux_C48_N30198_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C48_N30198_O_3_C_6_io_config = configBlock_ioBundle_confOut[622:619]; // @[TileFull.scala 151:60]
  assign SBMux_C48_N30198_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C48_N30198_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C48_N30198_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C48_N30198_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C56_N30200_O_3_C_6_io_in = {SBMux_C56_N30200_O_3_C_6_io_in_hi,SBMux_C56_N30200_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C56_N30200_O_3_C_6_io_config = configBlock_ioBundle_confOut[626:623]; // @[TileFull.scala 151:60]
  assign SBMux_C56_N30200_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C56_N30200_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C56_N30200_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C56_N30200_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C64_N30202_O_3_C_7_io_in = {SBMux_C64_N30202_O_3_C_7_io_in_hi,SBMux_C64_N30202_O_3_C_7_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C64_N30202_O_3_C_7_io_config = configBlock_ioBundle_confOut[630:627]; // @[TileFull.scala 151:60]
  assign SBMux_C64_N30202_O_3_C_7_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C64_N30202_O_3_C_7_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C64_N30202_O_3_C_7_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C64_N30202_O_3_C_7_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C72_N30204_O_3_C_6_io_in = {SBMux_C72_N30204_O_3_C_6_io_in_hi,SBMux_C72_N30204_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C72_N30204_O_3_C_6_io_config = configBlock_ioBundle_confOut[634:631]; // @[TileFull.scala 151:60]
  assign SBMux_C72_N30204_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C72_N30204_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C72_N30204_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C72_N30204_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C80_N30206_O_3_C_6_io_in = {SBMux_C80_N30206_O_3_C_6_io_in_hi,SBMux_C80_N30206_O_3_C_6_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C80_N30206_O_3_C_6_io_config = configBlock_ioBundle_confOut[638:635]; // @[TileFull.scala 151:60]
  assign SBMux_C80_N30206_O_3_C_6_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C80_N30206_O_3_C_6_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C80_N30206_O_3_C_6_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C80_N30206_O_3_C_6_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C88_N30208_O_4_C_5_io_in = {SBMux_C88_N30208_O_4_C_5_io_in_hi,SBMux_C88_N30208_O_4_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C88_N30208_O_4_C_5_io_config = configBlock_ioBundle_confOut[642:639]; // @[TileFull.scala 151:60]
  assign SBMux_C88_N30208_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C88_N30208_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C88_N30208_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C88_N30208_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C96_N30210_O_4_C_5_io_in = {SBMux_C96_N30210_O_4_C_5_io_in_hi,SBMux_C96_N30210_O_4_C_5_io_in_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C96_N30210_O_4_C_5_io_config = configBlock_ioBundle_confOut[646:643]; // @[TileFull.scala 151:60]
  assign SBMux_C96_N30210_O_4_C_5_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C96_N30210_O_4_C_5_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C96_N30210_O_4_C_5_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C96_N30210_O_4_C_5_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C100_N30212_O_4_C_1_io_in = {SBMux_C100_N30212_O_4_C_1_io_in_hi,SBMux_C0_N30186_O_4_C_6_io_in_lo_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C100_N30212_O_4_C_1_io_config = configBlock_ioBundle_confOut[649:647]; // @[TileFull.scala 151:60]
  assign SBMux_C100_N30212_O_4_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C100_N30212_O_4_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C100_N30212_O_4_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C100_N30212_O_4_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
  assign SBMux_C104_N30214_O_3_C_1_io_in = {SBMux_C104_N30214_O_3_C_1_io_in_hi,SBMux_C40_N30196_O_3_C_5_io_in_lo_lo}; // @[TileFull.scala 202:13]
  assign SBMux_C104_N30214_O_3_C_1_io_config = configBlock_ioBundle_confOut[652:650]; // @[TileFull.scala 151:60]
  assign SBMux_C104_N30214_O_3_C_1_io_loopBreak = ctrlSignals_loopBreak; // @[TileFull.scala 155:28]
  assign SBMux_C104_N30214_O_3_C_1_io_ioGndBle = ctrlSignals_gndBlkOuts; // @[TileFull.scala 158:27]
  assign SBMux_C104_N30214_O_3_C_1_io_cnstClk = ctrlSignals_constClock; // @[TileFull.scala 156:26]
  assign SBMux_C104_N30214_O_3_C_1_io_arst = ctrlSignals_arst; // @[TileFull.scala 157:23]
endmodule
